magic
tech scmos
timestamp 1590329367
<< metal1 >>
rect -2 97 34 103
rect 2 57 6 94
rect 10 60 14 94
rect 18 57 22 94
rect 2 54 22 57
rect 26 54 30 94
rect 26 50 29 54
rect 2 43 6 47
rect 9 44 10 49
rect 18 44 23 47
rect 10 40 14 41
rect 10 33 14 37
rect 18 26 21 44
rect 26 43 30 47
rect 5 6 9 26
rect 18 6 22 26
rect 26 23 30 27
rect 25 19 29 20
rect 26 6 30 16
rect -2 -3 34 3
<< labels >>
rlabel metal1 2 43 6 47 6 A
port 1 nsew default input
rlabel metal1 10 33 14 37 6 B
port 2 nsew default input
rlabel metal1 26 23 30 27 6 C
port 3 nsew default input
rlabel metal1 -2 -3 34 3 8 gnd
port 4 nsew ground bidirectional
rlabel metal1 26 43 30 47 6 Y
port 5 nsew default output
rlabel metal1 -2 97 34 103 6 vdd
port 6 nsew power bidirectional
<< properties >>
string LEFclass CORE
string LEFsite core
string LEFview TRUE
string FIXED_BBOX 0 0 32 100
string LEFsymmetry X Y
<< end >>
