magic
tech scmos
timestamp 1590329367
<< metal1 >>
rect -2 97 42 103
rect 2 54 6 94
rect 10 51 14 94
rect 18 54 22 94
rect 26 51 30 94
rect 34 54 38 94
rect 10 50 30 51
rect 10 47 23 50
rect 26 43 30 47
rect 2 33 6 37
rect 26 33 30 40
rect 2 29 6 30
rect 10 29 30 33
rect 2 6 6 26
rect 10 6 14 29
rect 18 6 22 26
rect 26 6 30 29
rect 34 6 38 26
rect -2 -3 42 3
<< labels >>
rlabel metal1 2 33 6 37 6 A
port 1 nsew default input
rlabel metal1 -2 -3 42 3 8 gnd
port 2 nsew ground bidirectional
rlabel metal1 26 43 30 47 6 Y
port 3 nsew default output
rlabel metal1 -2 97 42 103 6 vdd
port 4 nsew power bidirectional
<< properties >>
string LEFclass CORE
string LEFsite core
string LEFview TRUE
string FIXED_BBOX 0 0 40 100
string LEFsymmetry X Y
<< end >>
