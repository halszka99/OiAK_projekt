magic
tech scmos
timestamp 1590329367
<< metal1 >>
rect -2 97 34 103
rect 2 57 6 94
rect 10 60 14 94
rect 18 59 22 94
rect 2 54 15 57
rect 18 54 23 59
rect 26 54 30 94
rect 2 43 6 47
rect 12 44 15 54
rect 12 40 17 44
rect 20 40 23 54
rect 3 39 7 40
rect 12 32 15 40
rect 18 33 22 37
rect 2 29 15 32
rect 2 6 6 29
rect 20 26 23 30
rect 10 6 14 26
rect 18 23 23 26
rect 18 6 22 23
rect 26 6 30 26
rect -2 -3 34 3
<< labels >>
rlabel metal1 2 43 6 47 6 A
port 1 nsew default input
rlabel metal1 -2 -3 34 3 8 gnd
port 2 nsew ground bidirectional
rlabel metal1 18 33 22 37 6 Y
port 3 nsew default output
rlabel metal1 -2 97 34 103 6 vdd
port 4 nsew power bidirectional
<< properties >>
string LEFclass CORE
string LEFsite core
string LEFview TRUE
string FIXED_BBOX 0 0 32 100
string LEFsymmetry X Y
<< end >>
