magic
tech scmos
timestamp 1590329367
<< metal1 >>
rect -2 97 42 103
rect 2 54 6 94
rect 15 54 25 94
rect 34 54 38 94
rect 10 43 14 47
rect 18 40 21 54
rect 26 43 30 47
rect 34 40 38 41
rect 10 39 14 40
rect 26 39 30 40
rect 2 33 6 37
rect 9 31 10 36
rect 18 33 22 37
rect 25 33 30 36
rect 34 33 38 37
rect 3 26 21 28
rect 27 26 30 33
rect 2 25 22 26
rect 2 6 6 25
rect 10 6 14 22
rect 18 9 22 25
rect 26 12 30 26
rect 34 9 38 26
rect 18 6 38 9
rect -2 -3 42 3
<< labels >>
rlabel metal1 2 33 6 37 6 A
port 1 nsew default input
rlabel metal1 10 43 14 47 6 B
port 2 nsew default input
rlabel metal1 34 33 38 37 6 C
port 3 nsew default input
rlabel metal1 26 43 30 47 6 D
port 4 nsew default input
rlabel metal1 -2 -3 42 3 8 gnd
port 5 nsew ground bidirectional
rlabel metal1 18 33 22 37 6 Y
port 6 nsew default output
rlabel metal1 -2 97 42 103 6 vdd
port 7 nsew power bidirectional
<< properties >>
string LEFclass CORE
string LEFsite core
string LEFview TRUE
string FIXED_BBOX 0 0 40 100
string LEFsymmetry X Y
<< end >>
