VERSION 5.3 ;
   NAMESCASESENSITIVE ON ;
   NOWIREEXTENSIONATPIN ON ;
   DIVIDERCHAR "/" ;
   BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO in
   CLASS BLOCK ;
   FOREIGN in ;
   ORIGIN 3.3000 -0.6000 ;
   SIZE 85.6500 BY 42.3000 ;
   PIN x
      PORT
         LAYER metal1 ;
	    RECT 45.0000 24.4500 46.2000 24.6000 ;
	    RECT 45.0000 23.5500 53.2500 24.4500 ;
	    RECT 45.0000 23.4000 46.2000 23.5500 ;
	    RECT 52.3500 21.4500 53.2500 23.5500 ;
	    RECT 54.6000 21.4500 55.8000 21.6000 ;
	    RECT 52.3500 20.5500 55.8000 21.4500 ;
	    RECT 54.6000 20.4000 55.8000 20.5500 ;
         LAYER metal2 ;
	    RECT 42.6000 41.4000 43.8000 42.6000 ;
	    RECT 47.4000 41.4000 48.6000 42.6000 ;
	    RECT 42.7500 27.4500 43.6500 41.4000 ;
	    RECT 47.5500 35.5500 48.4500 41.4000 ;
	    RECT 42.7500 26.5500 46.0500 27.4500 ;
	    RECT 45.1500 24.6000 46.0500 26.5500 ;
	    RECT 45.0000 23.4000 46.2000 24.6000 ;
         LAYER metal3 ;
	    RECT 42.3000 42.7500 44.1000 42.9000 ;
	    RECT 47.1000 42.7500 48.9000 42.9000 ;
	    RECT 42.3000 41.2500 48.9000 42.7500 ;
	    RECT 42.3000 41.1000 44.1000 41.2500 ;
	    RECT 47.1000 41.1000 48.9000 41.2500 ;
      END
   END x
   PIN y
      PORT
         LAYER metal1 ;
	    RECT 40.2000 23.4000 41.4000 24.6000 ;
	    RECT 69.0000 20.4000 70.2000 21.6000 ;
         LAYER metal2 ;
	    RECT 40.3500 24.6000 41.2500 36.4500 ;
	    RECT 40.2000 23.4000 41.4000 24.6000 ;
	    RECT 69.0000 23.4000 70.2000 24.6000 ;
	    RECT 69.1500 21.6000 70.0500 23.4000 ;
	    RECT 69.0000 20.4000 70.2000 21.6000 ;
         LAYER metal3 ;
	    RECT 39.9000 24.7500 41.7000 24.9000 ;
	    RECT 68.7000 24.7500 70.5000 24.9000 ;
	    RECT 39.9000 23.2500 70.5000 24.7500 ;
	    RECT 39.9000 23.1000 41.7000 23.2500 ;
	    RECT 68.7000 23.1000 70.5000 23.2500 ;
      END
   END y
   PIN g
      PORT
         LAYER metal1 ;
	    RECT 9.0000 20.4000 10.2000 21.6000 ;
         LAYER metal2 ;
	    RECT -3.0000 36.4500 -1.8000 36.6000 ;
	    RECT -3.0000 35.5500 2.8500 36.4500 ;
	    RECT -3.0000 35.4000 -1.8000 35.5500 ;
	    RECT 1.9500 30.6000 2.8500 35.5500 ;
	    RECT 1.8000 29.4000 3.0000 30.6000 ;
	    RECT 9.0000 29.4000 10.2000 30.6000 ;
	    RECT 9.1500 21.6000 10.0500 29.4000 ;
	    RECT 9.0000 20.4000 10.2000 21.6000 ;
         LAYER metal3 ;
	    RECT -3.3000 35.1000 -1.5000 36.9000 ;
	    RECT -3.1500 29.2500 -1.6500 35.1000 ;
	    RECT 1.5000 30.7500 3.3000 30.9000 ;
	    RECT 8.7000 30.7500 10.5000 30.9000 ;
	    RECT 1.5000 29.2500 10.5000 30.7500 ;
	    RECT 1.5000 29.1000 3.3000 29.2500 ;
	    RECT 8.7000 29.1000 10.5000 29.2500 ;
      END
   END g
   PIN p
      PORT
         LAYER metal1 ;
	    RECT 1.8000 20.4000 3.0000 21.6000 ;
         LAYER metal2 ;
	    RECT 1.8000 20.4000 3.0000 21.6000 ;
	    RECT 1.9500 18.6000 2.8500 20.4000 ;
	    RECT 1.8000 17.4000 3.0000 18.6000 ;
         LAYER metal3 ;
	    RECT -3.1500 18.7500 -1.6500 24.7500 ;
	    RECT 1.5000 18.7500 3.3000 18.9000 ;
	    RECT -3.1500 17.2500 3.3000 18.7500 ;
	    RECT 1.5000 17.1000 3.3000 17.2500 ;
      END
   END p
   PIN h
      PORT
         LAYER metal1 ;
	    RECT 76.2000 20.4000 77.4000 21.6000 ;
         LAYER metal2 ;
	    RECT 76.2000 20.4000 77.4000 21.6000 ;
	    RECT 76.3500 18.6000 77.2500 20.4000 ;
	    RECT 76.2000 17.4000 77.4000 18.6000 ;
         LAYER metal3 ;
	    RECT 75.9000 18.7500 77.7000 18.9000 ;
	    RECT 80.8500 18.7500 82.3500 24.7500 ;
	    RECT 75.9000 17.2500 82.3500 18.7500 ;
	    RECT 75.9000 17.1000 77.7000 17.2500 ;
      END
   END h
   OBS
         LAYER metal1 ;
	    RECT 0.6000 30.6000 78.6000 32.4000 ;
	    RECT 1.8000 22.5000 3.0000 29.7000 ;
	    RECT 4.2000 23.7000 5.4000 29.7000 ;
	    RECT 6.6000 22.8000 7.8000 29.7000 ;
	    RECT 4.5000 21.9000 7.8000 22.8000 ;
	    RECT 9.0000 22.5000 10.2000 29.7000 ;
	    RECT 11.4000 23.7000 12.6000 29.7000 ;
	    RECT 13.8000 22.8000 15.0000 29.7000 ;
	    RECT 24.3000 24.6000 25.5000 29.7000 ;
	    RECT 24.3000 23.7000 27.0000 24.6000 ;
	    RECT 28.2000 23.7000 29.4000 29.7000 ;
	    RECT 30.6000 26.7000 31.8000 29.7000 ;
	    RECT 33.0000 26.7000 34.2000 29.7000 ;
	    RECT 35.4000 26.7000 36.6000 29.7000 ;
	    RECT 11.7000 21.9000 15.0000 22.8000 ;
	    RECT 1.8000 18.6000 3.0000 19.5000 ;
	    RECT 1.8000 15.3000 2.7000 18.6000 ;
	    RECT 4.5000 17.4000 5.4000 21.9000 ;
	    RECT 6.6000 19.5000 7.8000 19.8000 ;
	    RECT 9.0000 18.6000 10.2000 19.5000 ;
	    RECT 6.6000 17.4000 7.8000 18.6000 ;
	    RECT 3.6000 16.2000 5.4000 17.4000 ;
	    RECT 4.5000 15.3000 5.4000 16.2000 ;
	    RECT 9.0000 15.3000 9.9000 18.6000 ;
	    RECT 11.7000 17.4000 12.6000 21.9000 ;
	    RECT 18.6000 21.4500 19.8000 21.6000 ;
	    RECT 18.6000 20.5500 24.4500 21.4500 ;
	    RECT 18.6000 20.4000 19.8000 20.5500 ;
	    RECT 13.8000 19.5000 15.0000 19.8000 ;
	    RECT 13.8000 18.4500 15.0000 18.6000 ;
	    RECT 21.0000 18.4500 22.2000 18.6000 ;
	    RECT 13.8000 17.5500 22.2000 18.4500 ;
	    RECT 23.5500 18.4500 24.4500 20.5500 ;
	    RECT 25.8000 19.5000 27.0000 23.7000 ;
	    RECT 28.2000 22.5000 29.4000 22.8000 ;
	    RECT 33.0000 22.5000 33.9000 26.7000 ;
	    RECT 35.4000 25.5000 36.6000 25.8000 ;
	    RECT 35.4000 23.4000 36.6000 24.6000 ;
	    RECT 28.2000 20.4000 29.4000 21.6000 ;
	    RECT 30.6000 21.4500 31.8000 21.6000 ;
	    RECT 33.0000 21.4500 34.2000 21.6000 ;
	    RECT 30.6000 20.5500 34.2000 21.4500 ;
	    RECT 35.5500 21.4500 36.4500 23.4000 ;
	    RECT 37.8000 22.5000 39.0000 29.7000 ;
	    RECT 40.2000 26.7000 41.4000 29.7000 ;
	    RECT 40.2000 25.5000 41.4000 25.8000 ;
	    RECT 42.6000 22.5000 43.8000 29.7000 ;
	    RECT 45.0000 26.7000 46.2000 29.7000 ;
	    RECT 45.0000 25.5000 46.2000 25.8000 ;
	    RECT 54.6000 23.7000 55.8000 29.7000 ;
	    RECT 57.0000 24.6000 58.5000 29.7000 ;
	    RECT 61.2000 24.3000 63.6000 29.7000 ;
	    RECT 66.3000 24.6000 67.8000 29.7000 ;
	    RECT 54.6000 22.8000 58.2000 23.7000 ;
	    RECT 57.0000 22.5000 58.2000 22.8000 ;
	    RECT 59.1000 22.2000 60.3000 23.4000 ;
	    RECT 59.1000 21.6000 60.0000 22.2000 ;
	    RECT 37.8000 21.4500 39.0000 21.6000 ;
	    RECT 35.5500 20.5500 39.0000 21.4500 ;
	    RECT 30.6000 20.4000 31.8000 20.5500 ;
	    RECT 33.0000 20.4000 34.2000 20.5500 ;
	    RECT 37.8000 20.4000 39.0000 20.5500 ;
	    RECT 40.2000 21.4500 41.4000 21.6000 ;
	    RECT 42.6000 21.4500 43.8000 21.6000 ;
	    RECT 40.2000 20.5500 43.8000 21.4500 ;
	    RECT 40.2000 20.4000 41.4000 20.5500 ;
	    RECT 42.6000 20.4000 43.8000 20.5500 ;
	    RECT 56.7000 20.4000 57.0000 21.6000 ;
	    RECT 58.8000 20.4000 60.0000 21.6000 ;
	    RECT 61.2000 21.3000 62.1000 24.3000 ;
	    RECT 69.0000 23.7000 70.2000 29.7000 ;
	    RECT 63.0000 22.2000 65.4000 23.4000 ;
	    RECT 66.3000 22.8000 70.2000 23.7000 ;
	    RECT 71.4000 22.8000 72.6000 29.7000 ;
	    RECT 73.8000 23.7000 75.0000 29.7000 ;
	    RECT 66.3000 22.5000 67.5000 22.8000 ;
	    RECT 71.4000 21.9000 74.7000 22.8000 ;
	    RECT 76.2000 22.5000 77.4000 29.7000 ;
	    RECT 67.8000 21.3000 68.1000 21.6000 ;
	    RECT 61.2000 20.4000 62.7000 21.3000 ;
	    RECT 66.9000 21.0000 68.1000 21.3000 ;
	    RECT 61.8000 19.5000 62.7000 20.4000 ;
	    RECT 63.6000 20.4000 68.1000 21.0000 ;
	    RECT 63.6000 20.1000 67.8000 20.4000 ;
	    RECT 63.6000 19.8000 64.8000 20.1000 ;
	    RECT 71.4000 19.5000 72.6000 19.8000 ;
	    RECT 25.8000 18.4500 27.0000 18.6000 ;
	    RECT 23.5500 17.5500 27.0000 18.4500 ;
	    RECT 13.8000 17.4000 15.0000 17.5500 ;
	    RECT 21.0000 17.4000 22.2000 17.5500 ;
	    RECT 25.8000 17.4000 27.0000 17.5500 ;
	    RECT 30.6000 17.4000 31.8000 18.6000 ;
	    RECT 10.8000 16.2000 12.6000 17.4000 ;
	    RECT 11.7000 15.3000 12.6000 16.2000 ;
	    RECT 1.8000 3.3000 3.0000 15.3000 ;
	    RECT 4.5000 14.4000 7.8000 15.3000 ;
	    RECT 4.2000 3.3000 5.4000 13.5000 ;
	    RECT 6.6000 3.3000 7.8000 14.4000 ;
	    RECT 9.0000 3.3000 10.2000 15.3000 ;
	    RECT 11.7000 14.4000 15.0000 15.3000 ;
	    RECT 23.4000 14.4000 24.6000 15.6000 ;
	    RECT 11.4000 3.3000 12.6000 13.5000 ;
	    RECT 13.8000 3.3000 15.0000 14.4000 ;
	    RECT 23.4000 13.2000 24.6000 13.5000 ;
	    RECT 23.4000 3.3000 24.6000 9.3000 ;
	    RECT 25.8000 3.3000 27.0000 16.5000 ;
	    RECT 30.6000 16.2000 31.8000 16.5000 ;
	    RECT 33.0000 15.3000 33.9000 19.5000 ;
	    RECT 31.5000 14.1000 34.2000 15.3000 ;
	    RECT 28.2000 3.3000 29.4000 9.3000 ;
	    RECT 31.5000 3.3000 32.7000 14.1000 ;
	    RECT 35.4000 3.3000 36.6000 15.3000 ;
	    RECT 37.8000 3.3000 39.0000 19.5000 ;
	    RECT 40.2000 3.3000 41.4000 9.3000 ;
	    RECT 42.6000 3.3000 43.8000 19.5000 ;
	    RECT 61.8000 17.4000 63.0000 18.6000 ;
	    RECT 65.7000 18.3000 66.9000 18.6000 ;
	    RECT 64.5000 17.4000 66.9000 18.3000 ;
	    RECT 69.0000 18.4500 70.2000 18.6000 ;
	    RECT 71.4000 18.4500 72.6000 18.6000 ;
	    RECT 69.0000 17.5500 72.6000 18.4500 ;
	    RECT 69.0000 17.4000 70.2000 17.5500 ;
	    RECT 71.4000 17.4000 72.6000 17.5500 ;
	    RECT 73.8000 17.4000 74.7000 21.9000 ;
	    RECT 76.2000 18.6000 77.4000 19.5000 ;
	    RECT 64.5000 17.1000 65.7000 17.4000 ;
	    RECT 61.8000 15.3000 62.7000 16.5000 ;
	    RECT 73.8000 16.2000 75.6000 17.4000 ;
	    RECT 73.8000 15.3000 74.7000 16.2000 ;
	    RECT 76.5000 15.3000 77.4000 18.6000 ;
	    RECT 54.6000 14.4000 58.2000 15.3000 ;
	    RECT 45.0000 3.3000 46.2000 9.3000 ;
	    RECT 54.6000 3.3000 55.8000 14.4000 ;
	    RECT 57.0000 14.1000 58.2000 14.4000 ;
	    RECT 57.0000 3.3000 58.5000 13.2000 ;
	    RECT 61.2000 3.3000 63.6000 15.3000 ;
	    RECT 66.3000 14.4000 70.2000 15.3000 ;
	    RECT 66.3000 14.1000 67.5000 14.4000 ;
	    RECT 66.3000 3.3000 67.8000 13.2000 ;
	    RECT 69.0000 3.3000 70.2000 14.4000 ;
	    RECT 71.4000 14.4000 74.7000 15.3000 ;
	    RECT 71.4000 3.3000 72.6000 14.4000 ;
	    RECT 73.8000 3.3000 75.0000 13.5000 ;
	    RECT 76.2000 3.3000 77.4000 15.3000 ;
	    RECT 0.6000 0.6000 78.6000 2.4000 ;
         LAYER metal2 ;
	    RECT 46.8000 30.6000 54.0000 32.4000 ;
	    RECT 21.1500 26.5500 31.6500 27.4500 ;
	    RECT 18.6000 20.4000 19.8000 21.6000 ;
	    RECT 18.7500 18.6000 19.6500 20.4000 ;
	    RECT 21.1500 18.6000 22.0500 26.5500 ;
	    RECT 28.2000 23.4000 29.4000 24.6000 ;
	    RECT 28.3500 21.6000 29.2500 23.4000 ;
	    RECT 30.7500 21.6000 31.6500 26.5500 ;
	    RECT 35.4000 23.4000 36.6000 24.6000 ;
	    RECT 57.0000 22.5000 58.2000 23.7000 ;
	    RECT 66.3000 23.4000 67.5000 23.7000 ;
	    RECT 59.1000 22.5000 67.5000 23.4000 ;
	    RECT 28.2000 20.4000 29.4000 21.6000 ;
	    RECT 30.6000 20.4000 31.8000 21.6000 ;
	    RECT 40.2000 20.4000 41.4000 21.6000 ;
	    RECT 57.0000 21.3000 57.9000 22.5000 ;
	    RECT 59.1000 22.2000 60.3000 22.5000 ;
	    RECT 64.2000 22.2000 65.4000 22.5000 ;
	    RECT 57.0000 20.4000 65.4000 21.3000 ;
	    RECT 40.3500 18.6000 41.2500 20.4000 ;
	    RECT 6.6000 17.4000 7.8000 18.6000 ;
	    RECT 18.6000 17.4000 19.8000 18.6000 ;
	    RECT 21.0000 17.4000 22.2000 18.6000 ;
	    RECT 23.4000 17.4000 24.6000 18.6000 ;
	    RECT 30.6000 17.4000 31.8000 18.6000 ;
	    RECT 40.2000 17.4000 41.4000 18.6000 ;
	    RECT 23.5500 15.6000 24.4500 17.4000 ;
	    RECT 23.4000 14.4000 24.6000 15.6000 ;
	    RECT 57.0000 15.3000 57.9000 20.4000 ;
	    RECT 61.8000 17.4000 63.0000 18.6000 ;
	    RECT 64.5000 18.3000 65.4000 20.4000 ;
	    RECT 64.5000 17.1000 65.7000 18.3000 ;
	    RECT 66.6000 15.3000 67.5000 22.5000 ;
	    RECT 69.0000 17.4000 70.2000 18.6000 ;
	    RECT 57.0000 14.1000 58.2000 15.3000 ;
	    RECT 66.3000 14.1000 67.5000 15.3000 ;
	    RECT 15.6000 0.6000 22.8000 2.4000 ;
         LAYER metal3 ;
	    RECT 46.8000 30.6000 54.0000 32.4000 ;
	    RECT 27.9000 24.7500 29.7000 24.9000 ;
	    RECT 35.1000 24.7500 36.9000 24.9000 ;
	    RECT 27.9000 23.2500 36.9000 24.7500 ;
	    RECT 27.9000 23.1000 29.7000 23.2500 ;
	    RECT 35.1000 23.1000 36.9000 23.2500 ;
	    RECT 6.3000 18.7500 8.1000 18.9000 ;
	    RECT 18.3000 18.7500 20.1000 18.9000 ;
	    RECT 6.3000 17.2500 20.1000 18.7500 ;
	    RECT 6.3000 17.1000 8.1000 17.2500 ;
	    RECT 18.3000 17.1000 20.1000 17.2500 ;
	    RECT 23.1000 18.7500 24.9000 18.9000 ;
	    RECT 30.3000 18.7500 32.1000 18.9000 ;
	    RECT 39.9000 18.7500 41.7000 18.9000 ;
	    RECT 23.1000 17.2500 41.7000 18.7500 ;
	    RECT 23.1000 17.1000 24.9000 17.2500 ;
	    RECT 30.3000 17.1000 32.1000 17.2500 ;
	    RECT 39.9000 17.1000 41.7000 17.2500 ;
	    RECT 61.5000 18.7500 63.3000 18.9000 ;
	    RECT 68.7000 18.7500 70.5000 18.9000 ;
	    RECT 61.5000 17.2500 70.5000 18.7500 ;
	    RECT 61.5000 17.1000 63.3000 17.2500 ;
	    RECT 68.7000 17.1000 70.5000 17.2500 ;
	    RECT 15.6000 0.6000 22.8000 2.4000 ;
   END
END in
