* NGSPICE file created from dot.ext - technology: scmos

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

.subckt dot Gh Ph Gl Pl Ghl Phl
XNAND2X1_2 INVX1_1/Y NAND2X1_1/Y BUFX2_2/gnd BUFX2_1/A BUFX2_2/vdd NAND2X1
XFILL_0_0_2 BUFX2_2/gnd BUFX2_2/vdd FILL
XINVX1_1 Gh BUFX2_2/gnd INVX1_1/Y BUFX2_2/vdd INVX1
XAND2X2_1 Ph Pl BUFX2_2/gnd BUFX2_2/A BUFX2_2/vdd AND2X2
XFILL_0_1_0 BUFX2_2/gnd BUFX2_2/vdd FILL
XFILL_0_1_2 BUFX2_2/gnd BUFX2_2/vdd FILL
XFILL_0_1_1 BUFX2_2/gnd BUFX2_2/vdd FILL
XBUFX2_1 BUFX2_1/A BUFX2_2/gnd Ghl BUFX2_2/vdd BUFX2
XFILL_0_0_0 BUFX2_2/gnd BUFX2_2/vdd FILL
XNAND2X1_1 Gl Ph BUFX2_2/gnd NAND2X1_1/Y BUFX2_2/vdd NAND2X1
XFILL_0_0_1 BUFX2_2/gnd BUFX2_2/vdd FILL
XBUFX2_2 BUFX2_2/A BUFX2_2/gnd Phl BUFX2_2/vdd BUFX2
.ends

