VERSION 5.3 ;
   NAMESCASESENSITIVE ON ;
   NOWIREEXTENSIONATPIN ON ;
   DIVIDERCHAR "/" ;
   BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO adder
   CLASS BLOCK ;
   FOREIGN adder ;
   ORIGIN 3.1500 3.4500 ;
   SIZE 200.7000 BY 99.9000 ;
   PIN x0
      PORT
         LAYER metal1 ;
	    RECT 40.2000 83.4000 41.4000 84.6000 ;
	    RECT 23.4000 80.4000 24.6000 81.6000 ;
         LAYER metal2 ;
	    RECT 37.9500 95.5500 41.2500 96.4500 ;
	    RECT 40.3500 84.6000 41.2500 95.5500 ;
	    RECT 23.4000 83.4000 24.6000 84.6000 ;
	    RECT 40.2000 83.4000 41.4000 84.6000 ;
	    RECT 23.5500 81.6000 24.4500 83.4000 ;
	    RECT 23.4000 80.4000 24.6000 81.6000 ;
         LAYER metal3 ;
	    RECT 23.1000 84.7500 24.9000 84.9000 ;
	    RECT 39.9000 84.7500 41.7000 84.9000 ;
	    RECT 23.1000 83.2500 41.7000 84.7500 ;
	    RECT 23.1000 83.1000 24.9000 83.2500 ;
	    RECT 39.9000 83.1000 41.7000 83.2500 ;
      END
   END x0
   PIN x1
      PORT
         LAYER metal1 ;
	    RECT 109.8000 83.4000 111.0000 84.6000 ;
	    RECT 88.2000 80.4000 89.4000 81.6000 ;
         LAYER metal2 ;
	    RECT 109.9500 90.6000 110.8500 96.4500 ;
	    RECT 102.6000 89.4000 103.8000 90.6000 ;
	    RECT 109.8000 89.4000 111.0000 90.6000 ;
	    RECT 102.7500 87.4500 103.6500 89.4000 ;
	    RECT 100.3500 86.5500 103.6500 87.4500 ;
	    RECT 88.2000 83.4000 89.4000 84.6000 ;
	    RECT 95.4000 83.4000 96.6000 84.6000 ;
	    RECT 88.3500 81.6000 89.2500 83.4000 ;
	    RECT 88.2000 80.4000 89.4000 81.6000 ;
	    RECT 95.5500 81.4500 96.4500 83.4000 ;
	    RECT 100.3500 81.4500 101.2500 86.5500 ;
	    RECT 109.9500 84.6000 110.8500 89.4000 ;
	    RECT 109.8000 83.4000 111.0000 84.6000 ;
	    RECT 95.5500 80.5500 101.2500 81.4500 ;
         LAYER metal3 ;
	    RECT 102.3000 90.7500 104.1000 90.9000 ;
	    RECT 109.5000 90.7500 111.3000 90.9000 ;
	    RECT 102.3000 89.2500 111.3000 90.7500 ;
	    RECT 102.3000 89.1000 104.1000 89.2500 ;
	    RECT 109.5000 89.1000 111.3000 89.2500 ;
	    RECT 87.9000 84.7500 89.7000 84.9000 ;
	    RECT 95.1000 84.7500 96.9000 84.9000 ;
	    RECT 87.9000 83.2500 96.9000 84.7500 ;
	    RECT 87.9000 83.1000 89.7000 83.2500 ;
	    RECT 95.1000 83.1000 96.9000 83.2500 ;
      END
   END x1
   PIN x2
      PORT
         LAYER metal1 ;
	    RECT 157.8000 83.4000 159.0000 84.6000 ;
	    RECT 174.6000 80.4000 175.8000 81.6000 ;
         LAYER metal2 ;
	    RECT 153.1500 90.6000 154.0500 96.4500 ;
	    RECT 153.0000 89.4000 154.2000 90.6000 ;
	    RECT 157.8000 89.4000 159.0000 90.6000 ;
	    RECT 174.6000 89.4000 175.8000 90.6000 ;
	    RECT 157.9500 84.6000 158.8500 89.4000 ;
	    RECT 157.8000 83.4000 159.0000 84.6000 ;
	    RECT 174.7500 81.6000 175.6500 89.4000 ;
	    RECT 174.6000 80.4000 175.8000 81.6000 ;
         LAYER metal3 ;
	    RECT 152.7000 90.7500 154.5000 90.9000 ;
	    RECT 157.5000 90.7500 159.3000 90.9000 ;
	    RECT 174.3000 90.7500 176.1000 90.9000 ;
	    RECT 152.7000 89.2500 176.1000 90.7500 ;
	    RECT 152.7000 89.1000 154.5000 89.2500 ;
	    RECT 157.5000 89.1000 159.3000 89.2500 ;
	    RECT 174.3000 89.1000 176.1000 89.2500 ;
      END
   END x2
   PIN x3
      PORT
         LAYER metal1 ;
	    RECT 157.8000 23.4000 159.0000 24.6000 ;
	    RECT 179.4000 20.4000 180.6000 21.6000 ;
         LAYER metal2 ;
	    RECT 157.8000 23.4000 159.0000 24.6000 ;
	    RECT 157.9500 6.6000 158.8500 23.4000 ;
	    RECT 179.4000 20.4000 180.6000 21.6000 ;
	    RECT 179.5500 18.6000 180.4500 20.4000 ;
	    RECT 172.2000 17.4000 173.4000 18.6000 ;
	    RECT 179.4000 17.4000 180.6000 18.6000 ;
	    RECT 172.3500 6.6000 173.2500 17.4000 ;
	    RECT 157.8000 5.4000 159.0000 6.6000 ;
	    RECT 172.2000 5.4000 173.4000 6.6000 ;
	    RECT 172.3500 -3.4500 173.2500 5.4000 ;
         LAYER metal3 ;
	    RECT 171.9000 18.7500 173.7000 18.9000 ;
	    RECT 179.1000 18.7500 180.9000 18.9000 ;
	    RECT 171.9000 17.2500 180.9000 18.7500 ;
	    RECT 171.9000 17.1000 173.7000 17.2500 ;
	    RECT 179.1000 17.1000 180.9000 17.2500 ;
	    RECT 157.5000 6.7500 159.3000 6.9000 ;
	    RECT 171.9000 6.7500 173.7000 6.9000 ;
	    RECT 157.5000 5.2500 173.7000 6.7500 ;
	    RECT 157.5000 5.1000 159.3000 5.2500 ;
	    RECT 171.9000 5.1000 173.7000 5.2500 ;
      END
   END x3
   PIN x4
      PORT
         LAYER metal1 ;
	    RECT 90.6000 38.4000 91.8000 39.6000 ;
	    RECT 126.6000 20.4000 127.8000 21.6000 ;
	    RECT 121.8000 18.4500 123.0000 18.6000 ;
	    RECT 126.7500 18.4500 127.6500 20.4000 ;
	    RECT 121.8000 17.5500 127.6500 18.4500 ;
	    RECT 121.8000 17.4000 123.0000 17.5500 ;
         LAYER metal2 ;
	    RECT 90.6000 38.4000 91.8000 39.6000 ;
	    RECT 90.7500 12.6000 91.6500 38.4000 ;
	    RECT 121.8000 17.4000 123.0000 18.6000 ;
	    RECT 90.6000 11.4000 91.8000 12.6000 ;
	    RECT 119.4000 12.4500 120.6000 12.6000 ;
	    RECT 121.9500 12.4500 122.8500 17.4000 ;
	    RECT 119.4000 11.5500 122.8500 12.4500 ;
	    RECT 119.4000 11.4000 120.6000 11.5500 ;
	    RECT 119.5500 -3.4500 120.4500 11.4000 ;
         LAYER metal3 ;
	    RECT 90.3000 12.7500 92.1000 12.9000 ;
	    RECT 119.1000 12.7500 120.9000 12.9000 ;
	    RECT 90.3000 11.2500 120.9000 12.7500 ;
	    RECT 90.3000 11.1000 92.1000 11.2500 ;
	    RECT 119.1000 11.1000 120.9000 11.2500 ;
      END
   END x4
   PIN x5
      PORT
         LAYER metal1 ;
	    RECT 16.2000 41.4000 17.4000 42.6000 ;
	    RECT 6.6000 23.4000 7.8000 24.6000 ;
         LAYER metal2 ;
	    RECT 16.2000 41.4000 17.4000 42.6000 ;
	    RECT 16.3500 36.6000 17.2500 41.4000 ;
	    RECT 6.6000 35.4000 7.8000 36.6000 ;
	    RECT 16.2000 35.4000 17.4000 36.6000 ;
	    RECT 6.7500 30.6000 7.6500 35.4000 ;
	    RECT 6.6000 29.4000 7.8000 30.6000 ;
	    RECT 6.7500 24.6000 7.6500 29.4000 ;
	    RECT 6.6000 23.4000 7.8000 24.6000 ;
         LAYER metal3 ;
	    RECT 6.3000 36.7500 8.1000 36.9000 ;
	    RECT 15.9000 36.7500 17.7000 36.9000 ;
	    RECT 6.3000 35.2500 17.7000 36.7500 ;
	    RECT 6.3000 35.1000 8.1000 35.2500 ;
	    RECT 15.9000 35.1000 17.7000 35.2500 ;
	    RECT 6.3000 30.7500 8.1000 30.9000 ;
	    RECT -3.1500 29.2500 8.1000 30.7500 ;
	    RECT -3.1500 23.2500 -1.6500 29.2500 ;
	    RECT 6.3000 29.1000 8.1000 29.2500 ;
      END
   END x5
   PIN y0
      PORT
         LAYER metal1 ;
	    RECT 25.8000 83.4000 27.0000 84.6000 ;
	    RECT 9.0000 80.4000 10.2000 81.6000 ;
         LAYER metal2 ;
	    RECT 25.9500 90.6000 26.8500 96.4500 ;
	    RECT 9.0000 89.4000 10.2000 90.6000 ;
	    RECT 25.8000 89.4000 27.0000 90.6000 ;
	    RECT 9.1500 81.6000 10.0500 89.4000 ;
	    RECT 25.9500 84.6000 26.8500 89.4000 ;
	    RECT 25.8000 83.4000 27.0000 84.6000 ;
	    RECT 9.0000 80.4000 10.2000 81.6000 ;
         LAYER metal3 ;
	    RECT 8.7000 90.7500 10.5000 90.9000 ;
	    RECT 25.5000 90.7500 27.3000 90.9000 ;
	    RECT 8.7000 89.2500 27.3000 90.7500 ;
	    RECT 8.7000 89.1000 10.5000 89.2500 ;
	    RECT 25.5000 89.1000 27.3000 89.2500 ;
      END
   END y0
   PIN y1
      PORT
         LAYER metal1 ;
	    RECT 97.8000 83.4000 99.0000 84.6000 ;
	    RECT 73.8000 80.4000 75.0000 81.6000 ;
         LAYER metal2 ;
	    RECT 97.9500 90.6000 98.8500 96.4500 ;
	    RECT 73.8000 89.4000 75.0000 90.6000 ;
	    RECT 97.8000 89.4000 99.0000 90.6000 ;
	    RECT 73.9500 81.6000 74.8500 89.4000 ;
	    RECT 97.9500 84.6000 98.8500 89.4000 ;
	    RECT 97.8000 83.4000 99.0000 84.6000 ;
	    RECT 73.8000 80.4000 75.0000 81.6000 ;
         LAYER metal3 ;
	    RECT 73.5000 90.7500 75.3000 90.9000 ;
	    RECT 97.5000 90.7500 99.3000 90.9000 ;
	    RECT 73.5000 89.2500 99.3000 90.7500 ;
	    RECT 73.5000 89.1000 75.3000 89.2500 ;
	    RECT 97.5000 89.1000 99.3000 89.2500 ;
      END
   END y1
   PIN y2
      PORT
         LAYER metal1 ;
	    RECT 160.2000 80.4000 161.4000 81.6000 ;
	    RECT 165.0000 38.4000 166.2000 39.6000 ;
         LAYER metal2 ;
	    RECT 160.3500 95.5500 163.6500 96.4500 ;
	    RECT 160.3500 81.6000 161.2500 95.5500 ;
	    RECT 160.2000 80.4000 161.4000 81.6000 ;
	    RECT 160.3500 60.6000 161.2500 80.4000 ;
	    RECT 160.2000 59.4000 161.4000 60.6000 ;
	    RECT 165.0000 59.4000 166.2000 60.6000 ;
	    RECT 165.1500 39.6000 166.0500 59.4000 ;
	    RECT 165.0000 38.4000 166.2000 39.6000 ;
         LAYER metal3 ;
	    RECT 159.9000 60.7500 161.7000 60.9000 ;
	    RECT 164.7000 60.7500 166.5000 60.9000 ;
	    RECT 159.9000 59.2500 166.5000 60.7500 ;
	    RECT 159.9000 59.1000 161.7000 59.2500 ;
	    RECT 164.7000 59.1000 166.5000 59.2500 ;
      END
   END y2
   PIN y3
      PORT
         LAYER metal1 ;
	    RECT 162.6000 23.4000 163.8000 24.6000 ;
	    RECT 162.7500 21.6000 163.6500 23.4000 ;
	    RECT 162.6000 21.4500 163.8000 21.6000 ;
	    RECT 165.0000 21.4500 166.2000 21.6000 ;
	    RECT 162.6000 20.5500 166.2000 21.4500 ;
	    RECT 162.6000 20.4000 163.8000 20.5500 ;
	    RECT 165.0000 20.4000 166.2000 20.5500 ;
         LAYER metal2 ;
	    RECT 162.6000 20.4000 163.8000 21.6000 ;
	    RECT 162.7500 -2.5500 163.6500 20.4000 ;
	    RECT 160.3500 -3.4500 163.6500 -2.5500 ;
      END
   END y3
   PIN y4
      PORT
         LAYER metal1 ;
	    RECT 85.8000 38.4000 87.0000 39.6000 ;
	    RECT 112.2000 20.4000 113.4000 21.6000 ;
         LAYER metal2 ;
	    RECT 85.8000 38.4000 87.0000 39.6000 ;
	    RECT 85.9500 36.6000 86.8500 38.4000 ;
	    RECT 85.8000 35.4000 87.0000 36.6000 ;
	    RECT 93.0000 35.4000 94.2000 36.6000 ;
	    RECT 105.0000 35.4000 106.2000 36.6000 ;
	    RECT 93.1500 6.6000 94.0500 35.4000 ;
	    RECT 105.1500 30.6000 106.0500 35.4000 ;
	    RECT 105.0000 29.4000 106.2000 30.6000 ;
	    RECT 112.2000 29.4000 113.4000 30.6000 ;
	    RECT 112.3500 21.6000 113.2500 29.4000 ;
	    RECT 112.2000 20.4000 113.4000 21.6000 ;
	    RECT 93.0000 5.4000 94.2000 6.6000 ;
	    RECT 112.2000 5.4000 113.4000 6.6000 ;
	    RECT 112.3500 -3.4500 113.2500 5.4000 ;
         LAYER metal3 ;
	    RECT 85.5000 36.7500 87.3000 36.9000 ;
	    RECT 92.7000 36.7500 94.5000 36.9000 ;
	    RECT 104.7000 36.7500 106.5000 36.9000 ;
	    RECT 85.5000 35.2500 106.5000 36.7500 ;
	    RECT 85.5000 35.1000 87.3000 35.2500 ;
	    RECT 92.7000 35.1000 94.5000 35.2500 ;
	    RECT 104.7000 35.1000 106.5000 35.2500 ;
	    RECT 104.7000 30.7500 106.5000 30.9000 ;
	    RECT 111.9000 30.7500 113.7000 30.9000 ;
	    RECT 104.7000 29.2500 113.7000 30.7500 ;
	    RECT 104.7000 29.1000 106.5000 29.2500 ;
	    RECT 111.9000 29.1000 113.7000 29.2500 ;
	    RECT 92.7000 6.7500 94.5000 6.9000 ;
	    RECT 111.9000 6.7500 113.7000 6.9000 ;
	    RECT 92.7000 5.2500 113.7000 6.7500 ;
	    RECT 92.7000 5.1000 94.5000 5.2500 ;
	    RECT 111.9000 5.1000 113.7000 5.2500 ;
      END
   END y4
   PIN y5
      PORT
         LAYER metal1 ;
	    RECT 1.8000 41.4000 3.0000 42.6000 ;
	    RECT 1.8000 23.4000 3.0000 24.6000 ;
         LAYER metal2 ;
	    RECT 1.8000 41.4000 3.0000 42.6000 ;
	    RECT 1.9500 36.6000 2.8500 41.4000 ;
	    RECT 1.8000 35.4000 3.0000 36.6000 ;
	    RECT 1.9500 24.6000 2.8500 35.4000 ;
	    RECT 1.8000 23.4000 3.0000 24.6000 ;
         LAYER metal3 ;
	    RECT -3.1500 36.7500 -1.6500 42.7500 ;
	    RECT 1.5000 36.7500 3.3000 36.9000 ;
	    RECT -3.1500 35.2500 3.3000 36.7500 ;
	    RECT 1.5000 35.1000 3.3000 35.2500 ;
      END
   END y5
   PIN s0
      PORT
         LAYER metal1 ;
	    RECT 1.8000 80.4000 3.0000 81.6000 ;
         LAYER metal2 ;
	    RECT 1.8000 80.4000 3.0000 81.6000 ;
	    RECT 1.9500 78.6000 2.8500 80.4000 ;
	    RECT 1.8000 77.4000 3.0000 78.6000 ;
         LAYER metal3 ;
	    RECT 1.5000 78.7500 3.3000 78.9000 ;
	    RECT -3.1500 77.2500 3.3000 78.7500 ;
	    RECT -3.1500 71.2500 -1.6500 77.2500 ;
	    RECT 1.5000 77.1000 3.3000 77.2500 ;
      END
   END s0
   PIN s1
      PORT
         LAYER metal1 ;
	    RECT 42.6000 80.4000 43.8000 81.6000 ;
         LAYER metal2 ;
	    RECT 42.7500 95.5500 46.0500 96.4500 ;
	    RECT 42.7500 81.6000 43.6500 95.5500 ;
	    RECT 42.6000 80.4000 43.8000 81.6000 ;
      END
   END s1
   PIN s2
      PORT
         LAYER metal1 ;
	    RECT 186.6000 21.4500 187.8000 21.6000 ;
	    RECT 191.4000 21.4500 192.6000 21.6000 ;
	    RECT 186.6000 20.5500 192.6000 21.4500 ;
	    RECT 186.6000 20.4000 187.8000 20.5500 ;
	    RECT 191.4000 20.4000 192.6000 20.5500 ;
         LAYER metal2 ;
	    RECT 191.4000 20.4000 192.6000 21.6000 ;
	    RECT 191.5500 18.6000 192.4500 20.4000 ;
	    RECT 191.4000 17.4000 192.6000 18.6000 ;
         LAYER metal3 ;
	    RECT 191.1000 18.7500 192.9000 18.9000 ;
	    RECT 191.1000 17.2500 197.5500 18.7500 ;
	    RECT 191.1000 17.1000 192.9000 17.2500 ;
	    RECT 196.0500 11.2500 197.5500 17.2500 ;
      END
   END s2
   PIN s3
      PORT
         LAYER metal1 ;
	    RECT 189.0000 42.4500 190.2000 42.6000 ;
	    RECT 191.4000 42.4500 192.6000 42.6000 ;
	    RECT 189.0000 41.5500 192.6000 42.4500 ;
	    RECT 189.0000 41.4000 190.2000 41.5500 ;
	    RECT 191.4000 41.4000 192.6000 41.5500 ;
         LAYER metal2 ;
	    RECT 191.4000 47.4000 192.6000 48.6000 ;
	    RECT 191.5500 42.6000 192.4500 47.4000 ;
	    RECT 191.4000 41.4000 192.6000 42.6000 ;
         LAYER metal3 ;
	    RECT 191.1000 48.7500 192.9000 48.9000 ;
	    RECT 191.1000 47.2500 197.5500 48.7500 ;
	    RECT 191.1000 47.1000 192.9000 47.2500 ;
	    RECT 196.0500 41.2500 197.5500 47.2500 ;
      END
   END s3
   PIN s4
      PORT
         LAYER metal1 ;
	    RECT 88.2000 20.4000 89.4000 21.6000 ;
         LAYER metal2 ;
	    RECT 88.2000 20.4000 89.4000 21.6000 ;
	    RECT 88.3500 -2.5500 89.2500 20.4000 ;
	    RECT 88.3500 -3.4500 91.6500 -2.5500 ;
      END
   END s4
   PIN s5
      PORT
         LAYER metal1 ;
	    RECT 18.6000 41.4000 19.8000 42.6000 ;
         LAYER metal2 ;
	    RECT 18.6000 47.4000 19.8000 48.6000 ;
	    RECT 18.7500 42.6000 19.6500 47.4000 ;
	    RECT 18.6000 41.4000 19.8000 42.6000 ;
         LAYER metal3 ;
	    RECT -3.1500 48.7500 -1.6500 54.7500 ;
	    RECT 18.3000 48.7500 20.1000 48.9000 ;
	    RECT -3.1500 47.2500 20.1000 48.7500 ;
	    RECT 18.3000 47.1000 20.1000 47.2500 ;
      END
   END s5
   PIN ov
      PORT
         LAYER metal1 ;
	    RECT 85.8000 20.4000 87.0000 21.6000 ;
         LAYER metal2 ;
	    RECT 85.8000 20.4000 87.0000 21.6000 ;
	    RECT 85.9500 -2.5500 86.8500 20.4000 ;
	    RECT 83.5500 -3.4500 86.8500 -2.5500 ;
      END
   END ov
   OBS
         LAYER metal1 ;
	    RECT 0.6000 90.6000 193.8000 92.4000 ;
	    RECT 1.8000 82.5000 3.0000 89.7000 ;
	    RECT 4.2000 83.7000 5.4000 89.7000 ;
	    RECT 6.6000 82.8000 7.8000 89.7000 ;
	    RECT 9.0000 83.7000 10.2000 89.7000 ;
	    RECT 11.4000 84.6000 12.9000 89.7000 ;
	    RECT 15.6000 84.3000 18.0000 89.7000 ;
	    RECT 20.7000 84.6000 22.2000 89.7000 ;
	    RECT 9.0000 82.8000 12.9000 83.7000 ;
	    RECT 4.5000 81.9000 7.8000 82.8000 ;
	    RECT 11.7000 82.5000 12.9000 82.8000 ;
	    RECT 13.8000 82.2000 16.2000 83.4000 ;
	    RECT 1.8000 78.6000 3.0000 79.5000 ;
	    RECT 1.8000 75.3000 2.7000 78.6000 ;
	    RECT 4.5000 77.4000 5.4000 81.9000 ;
	    RECT 11.1000 81.3000 11.4000 81.6000 ;
	    RECT 17.1000 81.3000 18.0000 84.3000 ;
	    RECT 23.4000 83.7000 24.6000 89.7000 ;
	    RECT 25.8000 86.7000 27.0000 89.7000 ;
	    RECT 25.8000 85.5000 27.0000 85.8000 ;
	    RECT 18.9000 82.2000 20.1000 83.4000 ;
	    RECT 21.0000 82.8000 24.6000 83.7000 ;
	    RECT 21.0000 82.5000 22.2000 82.8000 ;
	    RECT 28.2000 82.5000 29.4000 89.7000 ;
	    RECT 30.6000 86.7000 31.8000 89.7000 ;
	    RECT 33.0000 86.7000 34.2000 89.7000 ;
	    RECT 35.4000 86.7000 36.6000 89.7000 ;
	    RECT 30.6000 85.5000 31.8000 85.8000 ;
	    RECT 30.6000 83.4000 31.8000 84.6000 ;
	    RECT 11.1000 81.0000 12.3000 81.3000 ;
	    RECT 11.1000 80.4000 15.6000 81.0000 ;
	    RECT 11.4000 80.1000 15.6000 80.4000 ;
	    RECT 14.4000 79.8000 15.6000 80.1000 ;
	    RECT 16.5000 80.4000 18.0000 81.3000 ;
	    RECT 19.2000 81.6000 20.1000 82.2000 ;
	    RECT 19.2000 80.4000 20.4000 81.6000 ;
	    RECT 22.2000 80.4000 22.5000 81.6000 ;
	    RECT 28.2000 81.4500 29.4000 81.6000 ;
	    RECT 30.7500 81.4500 31.6500 83.4000 ;
	    RECT 33.3000 82.5000 34.2000 86.7000 ;
	    RECT 37.8000 82.5000 39.0000 89.7000 ;
	    RECT 40.2000 86.7000 41.4000 89.7000 ;
	    RECT 40.2000 85.5000 41.4000 85.8000 ;
	    RECT 42.6000 82.5000 43.8000 89.7000 ;
	    RECT 45.0000 83.7000 46.2000 89.7000 ;
	    RECT 47.4000 82.8000 48.6000 89.7000 ;
	    RECT 57.0000 83.7000 58.2000 89.7000 ;
	    RECT 59.4000 84.6000 60.9000 89.7000 ;
	    RECT 63.6000 84.3000 66.0000 89.7000 ;
	    RECT 68.7000 84.6000 70.2000 89.7000 ;
	    RECT 57.0000 82.8000 60.6000 83.7000 ;
	    RECT 45.3000 81.9000 48.6000 82.8000 ;
	    RECT 59.4000 82.5000 60.6000 82.8000 ;
	    RECT 61.5000 82.2000 62.7000 83.4000 ;
	    RECT 28.2000 80.5500 31.6500 81.4500 ;
	    RECT 28.2000 80.4000 29.4000 80.5500 ;
	    RECT 33.0000 80.4000 34.2000 81.6000 ;
	    RECT 37.8000 81.4500 39.0000 81.6000 ;
	    RECT 35.5500 80.5500 39.0000 81.4500 ;
	    RECT 6.6000 79.5000 7.8000 79.8000 ;
	    RECT 16.5000 79.5000 17.4000 80.4000 ;
	    RECT 6.6000 78.4500 7.8000 78.6000 ;
	    RECT 9.0000 78.4500 10.2000 78.6000 ;
	    RECT 6.6000 77.5500 10.2000 78.4500 ;
	    RECT 6.6000 77.4000 7.8000 77.5500 ;
	    RECT 9.0000 77.4000 10.2000 77.5500 ;
	    RECT 12.3000 78.3000 13.5000 78.6000 ;
	    RECT 12.3000 77.4000 14.7000 78.3000 ;
	    RECT 16.2000 77.4000 17.4000 78.6000 ;
	    RECT 3.6000 76.2000 5.4000 77.4000 ;
	    RECT 13.5000 77.1000 14.7000 77.4000 ;
	    RECT 4.5000 75.3000 5.4000 76.2000 ;
	    RECT 16.5000 75.3000 17.4000 76.5000 ;
	    RECT 1.8000 63.3000 3.0000 75.3000 ;
	    RECT 4.5000 74.4000 7.8000 75.3000 ;
	    RECT 4.2000 63.3000 5.4000 73.5000 ;
	    RECT 6.6000 63.3000 7.8000 74.4000 ;
	    RECT 9.0000 74.4000 12.9000 75.3000 ;
	    RECT 9.0000 63.3000 10.2000 74.4000 ;
	    RECT 11.7000 74.1000 12.9000 74.4000 ;
	    RECT 11.4000 63.3000 12.9000 73.2000 ;
	    RECT 15.6000 63.3000 18.0000 75.3000 ;
	    RECT 21.0000 74.4000 24.6000 75.3000 ;
	    RECT 21.0000 74.1000 22.2000 74.4000 ;
	    RECT 20.7000 63.3000 22.2000 73.2000 ;
	    RECT 23.4000 63.3000 24.6000 74.4000 ;
	    RECT 25.8000 63.3000 27.0000 69.3000 ;
	    RECT 28.2000 63.3000 29.4000 79.5000 ;
	    RECT 33.3000 75.3000 34.2000 79.5000 ;
	    RECT 35.5500 78.6000 36.4500 80.5500 ;
	    RECT 37.8000 80.4000 39.0000 80.5500 ;
	    RECT 35.4000 77.4000 36.6000 78.6000 ;
	    RECT 35.4000 76.2000 36.6000 76.5000 ;
	    RECT 30.6000 63.3000 31.8000 75.3000 ;
	    RECT 33.0000 74.1000 35.7000 75.3000 ;
	    RECT 34.5000 63.3000 35.7000 74.1000 ;
	    RECT 37.8000 63.3000 39.0000 79.5000 ;
	    RECT 42.6000 78.6000 43.8000 79.5000 ;
	    RECT 42.6000 75.3000 43.5000 78.6000 ;
	    RECT 45.3000 77.4000 46.2000 81.9000 ;
	    RECT 61.5000 81.6000 62.4000 82.2000 ;
	    RECT 49.8000 81.4500 51.0000 81.6000 ;
	    RECT 57.0000 81.4500 58.2000 81.6000 ;
	    RECT 49.8000 80.5500 58.2000 81.4500 ;
	    RECT 49.8000 80.4000 51.0000 80.5500 ;
	    RECT 57.0000 80.4000 58.2000 80.5500 ;
	    RECT 59.1000 80.4000 59.4000 81.6000 ;
	    RECT 61.2000 80.4000 62.4000 81.6000 ;
	    RECT 63.6000 81.3000 64.5000 84.3000 ;
	    RECT 71.4000 83.7000 72.6000 89.7000 ;
	    RECT 65.4000 82.2000 67.8000 83.4000 ;
	    RECT 68.7000 82.8000 72.6000 83.7000 ;
	    RECT 73.8000 83.7000 75.0000 89.7000 ;
	    RECT 76.2000 84.6000 77.7000 89.7000 ;
	    RECT 80.4000 84.3000 82.8000 89.7000 ;
	    RECT 85.5000 84.6000 87.0000 89.7000 ;
	    RECT 73.8000 82.8000 77.7000 83.7000 ;
	    RECT 68.7000 82.5000 69.9000 82.8000 ;
	    RECT 76.5000 82.5000 77.7000 82.8000 ;
	    RECT 78.6000 82.2000 81.0000 83.4000 ;
	    RECT 70.2000 81.3000 70.5000 81.6000 ;
	    RECT 63.6000 80.4000 65.1000 81.3000 ;
	    RECT 69.3000 81.0000 70.5000 81.3000 ;
	    RECT 47.4000 79.5000 48.6000 79.8000 ;
	    RECT 64.2000 79.5000 65.1000 80.4000 ;
	    RECT 66.0000 80.4000 70.5000 81.0000 ;
	    RECT 71.4000 80.4000 72.6000 81.6000 ;
	    RECT 75.9000 81.3000 76.2000 81.6000 ;
	    RECT 81.9000 81.3000 82.8000 84.3000 ;
	    RECT 88.2000 83.7000 89.4000 89.7000 ;
	    RECT 90.6000 83.7000 91.8000 89.7000 ;
	    RECT 94.5000 84.6000 95.7000 89.7000 ;
	    RECT 97.8000 86.7000 99.0000 89.7000 ;
	    RECT 97.8000 85.5000 99.0000 85.8000 ;
	    RECT 93.0000 83.7000 95.7000 84.6000 ;
	    RECT 83.7000 82.2000 84.9000 83.4000 ;
	    RECT 85.8000 82.8000 89.4000 83.7000 ;
	    RECT 85.8000 82.5000 87.0000 82.8000 ;
	    RECT 90.6000 82.5000 91.8000 82.8000 ;
	    RECT 75.9000 81.0000 77.1000 81.3000 ;
	    RECT 75.9000 80.4000 80.4000 81.0000 ;
	    RECT 66.0000 80.1000 70.2000 80.4000 ;
	    RECT 76.2000 80.1000 80.4000 80.4000 ;
	    RECT 66.0000 79.8000 67.2000 80.1000 ;
	    RECT 79.2000 79.8000 80.4000 80.1000 ;
	    RECT 81.3000 80.4000 82.8000 81.3000 ;
	    RECT 84.0000 81.6000 84.9000 82.2000 ;
	    RECT 84.0000 80.4000 85.2000 81.6000 ;
	    RECT 87.0000 80.4000 87.3000 81.6000 ;
	    RECT 90.6000 80.4000 91.8000 81.6000 ;
	    RECT 81.3000 79.5000 82.2000 80.4000 ;
	    RECT 93.0000 79.5000 94.2000 83.7000 ;
	    RECT 100.2000 82.5000 101.4000 89.7000 ;
	    RECT 102.6000 83.7000 103.8000 89.7000 ;
	    RECT 106.5000 84.6000 107.7000 89.7000 ;
	    RECT 109.8000 86.7000 111.0000 89.7000 ;
	    RECT 109.8000 85.5000 111.0000 85.8000 ;
	    RECT 105.0000 83.7000 107.7000 84.6000 ;
	    RECT 102.6000 82.5000 103.8000 82.8000 ;
	    RECT 100.2000 81.4500 101.4000 81.6000 ;
	    RECT 102.6000 81.4500 103.8000 81.6000 ;
	    RECT 100.2000 80.5500 103.8000 81.4500 ;
	    RECT 100.2000 80.4000 101.4000 80.5500 ;
	    RECT 102.6000 80.4000 103.8000 80.5500 ;
	    RECT 105.0000 79.5000 106.2000 83.7000 ;
	    RECT 112.2000 82.5000 113.4000 89.7000 ;
	    RECT 114.6000 86.7000 115.8000 89.7000 ;
	    RECT 117.0000 86.7000 118.2000 89.7000 ;
	    RECT 119.4000 86.7000 120.6000 89.7000 ;
	    RECT 117.0000 82.5000 117.9000 86.7000 ;
	    RECT 119.4000 85.5000 120.6000 85.8000 ;
	    RECT 122.7000 84.6000 123.9000 89.7000 ;
	    RECT 119.4000 83.4000 120.6000 84.6000 ;
	    RECT 122.7000 83.7000 125.4000 84.6000 ;
	    RECT 126.6000 83.7000 127.8000 89.7000 ;
	    RECT 129.0000 86.7000 130.2000 89.7000 ;
	    RECT 129.0000 85.5000 130.2000 85.8000 ;
	    RECT 107.4000 81.4500 108.6000 81.6000 ;
	    RECT 112.2000 81.4500 113.4000 81.6000 ;
	    RECT 117.0000 81.4500 118.2000 81.6000 ;
	    RECT 121.8000 81.4500 123.0000 81.6000 ;
	    RECT 107.4000 80.5500 115.6500 81.4500 ;
	    RECT 107.4000 80.4000 108.6000 80.5500 ;
	    RECT 112.2000 80.4000 113.4000 80.5500 ;
	    RECT 47.4000 78.4500 48.6000 78.6000 ;
	    RECT 64.2000 78.4500 65.4000 78.6000 ;
	    RECT 47.4000 77.5500 65.4000 78.4500 ;
	    RECT 68.1000 78.3000 69.3000 78.6000 ;
	    RECT 47.4000 77.4000 48.6000 77.5500 ;
	    RECT 64.2000 77.4000 65.4000 77.5500 ;
	    RECT 66.9000 77.4000 69.3000 78.3000 ;
	    RECT 77.1000 78.3000 78.3000 78.6000 ;
	    RECT 77.1000 77.4000 79.5000 78.3000 ;
	    RECT 81.0000 77.4000 82.2000 78.6000 ;
	    RECT 93.0000 78.4500 94.2000 78.6000 ;
	    RECT 95.4000 78.4500 96.6000 78.6000 ;
	    RECT 93.0000 77.5500 96.6000 78.4500 ;
	    RECT 93.0000 77.4000 94.2000 77.5500 ;
	    RECT 95.4000 77.4000 96.6000 77.5500 ;
	    RECT 44.4000 76.2000 46.2000 77.4000 ;
	    RECT 66.9000 77.1000 68.1000 77.4000 ;
	    RECT 78.3000 77.1000 79.5000 77.4000 ;
	    RECT 45.3000 75.3000 46.2000 76.2000 ;
	    RECT 64.2000 75.3000 65.1000 76.5000 ;
	    RECT 81.3000 75.3000 82.2000 76.5000 ;
	    RECT 40.2000 63.3000 41.4000 69.3000 ;
	    RECT 42.6000 63.3000 43.8000 75.3000 ;
	    RECT 45.3000 74.4000 48.6000 75.3000 ;
	    RECT 45.0000 63.3000 46.2000 73.5000 ;
	    RECT 47.4000 63.3000 48.6000 74.4000 ;
	    RECT 57.0000 74.4000 60.6000 75.3000 ;
	    RECT 57.0000 63.3000 58.2000 74.4000 ;
	    RECT 59.4000 74.1000 60.6000 74.4000 ;
	    RECT 59.4000 63.3000 60.9000 73.2000 ;
	    RECT 63.6000 63.3000 66.0000 75.3000 ;
	    RECT 68.7000 74.4000 72.6000 75.3000 ;
	    RECT 68.7000 74.1000 69.9000 74.4000 ;
	    RECT 68.7000 63.3000 70.2000 73.2000 ;
	    RECT 71.4000 63.3000 72.6000 74.4000 ;
	    RECT 73.8000 74.4000 77.7000 75.3000 ;
	    RECT 73.8000 63.3000 75.0000 74.4000 ;
	    RECT 76.5000 74.1000 77.7000 74.4000 ;
	    RECT 76.2000 63.3000 77.7000 73.2000 ;
	    RECT 80.4000 63.3000 82.8000 75.3000 ;
	    RECT 85.8000 74.4000 89.4000 75.3000 ;
	    RECT 85.8000 74.1000 87.0000 74.4000 ;
	    RECT 85.5000 63.3000 87.0000 73.2000 ;
	    RECT 88.2000 63.3000 89.4000 74.4000 ;
	    RECT 90.6000 63.3000 91.8000 69.3000 ;
	    RECT 93.0000 63.3000 94.2000 76.5000 ;
	    RECT 95.4000 75.4500 96.6000 75.6000 ;
	    RECT 97.8000 75.4500 99.0000 75.6000 ;
	    RECT 95.4000 74.5500 99.0000 75.4500 ;
	    RECT 95.4000 74.4000 96.6000 74.5500 ;
	    RECT 97.8000 74.4000 99.0000 74.5500 ;
	    RECT 95.4000 73.2000 96.6000 73.5000 ;
	    RECT 95.4000 63.3000 96.6000 69.3000 ;
	    RECT 97.8000 63.3000 99.0000 69.3000 ;
	    RECT 100.2000 63.3000 101.4000 79.5000 ;
	    RECT 105.0000 77.4000 106.2000 78.6000 ;
	    RECT 102.6000 63.3000 103.8000 69.3000 ;
	    RECT 105.0000 63.3000 106.2000 76.5000 ;
	    RECT 107.4000 74.4000 108.6000 75.6000 ;
	    RECT 107.4000 73.2000 108.6000 73.5000 ;
	    RECT 107.4000 63.3000 108.6000 69.3000 ;
	    RECT 109.8000 63.3000 111.0000 69.3000 ;
	    RECT 112.2000 63.3000 113.4000 79.5000 ;
	    RECT 114.7500 78.6000 115.6500 80.5500 ;
	    RECT 117.0000 80.5500 123.0000 81.4500 ;
	    RECT 117.0000 80.4000 118.2000 80.5500 ;
	    RECT 121.8000 80.4000 123.0000 80.5500 ;
	    RECT 124.2000 79.5000 125.4000 83.7000 ;
	    RECT 129.0000 83.4000 130.2000 84.6000 ;
	    RECT 126.6000 82.5000 127.8000 82.8000 ;
	    RECT 131.4000 82.5000 132.6000 89.7000 ;
	    RECT 141.0000 83.7000 142.2000 89.7000 ;
	    RECT 144.9000 84.6000 146.1000 89.7000 ;
	    RECT 148.2000 86.7000 149.4000 89.7000 ;
	    RECT 150.6000 86.7000 151.8000 89.7000 ;
	    RECT 153.0000 86.7000 154.2000 89.7000 ;
	    RECT 143.4000 83.7000 146.1000 84.6000 ;
	    RECT 141.0000 82.5000 142.2000 82.8000 ;
	    RECT 126.6000 81.4500 127.8000 81.6000 ;
	    RECT 131.4000 81.4500 132.6000 81.6000 ;
	    RECT 126.6000 80.5500 132.6000 81.4500 ;
	    RECT 126.6000 80.4000 127.8000 80.5500 ;
	    RECT 131.4000 80.4000 132.6000 80.5500 ;
	    RECT 141.0000 80.4000 142.2000 81.6000 ;
	    RECT 143.4000 79.5000 144.6000 83.7000 ;
	    RECT 150.6000 82.5000 151.5000 86.7000 ;
	    RECT 153.0000 85.5000 154.2000 85.8000 ;
	    RECT 153.0000 83.4000 154.2000 84.6000 ;
	    RECT 155.4000 82.5000 156.6000 89.7000 ;
	    RECT 157.8000 86.7000 159.0000 89.7000 ;
	    RECT 157.8000 85.5000 159.0000 85.8000 ;
	    RECT 160.2000 83.7000 161.4000 89.7000 ;
	    RECT 162.6000 84.6000 164.1000 89.7000 ;
	    RECT 166.8000 84.3000 169.2000 89.7000 ;
	    RECT 171.9000 84.6000 173.4000 89.7000 ;
	    RECT 160.2000 82.8000 164.1000 83.7000 ;
	    RECT 162.9000 82.5000 164.1000 82.8000 ;
	    RECT 165.0000 82.2000 167.4000 83.4000 ;
	    RECT 145.8000 81.4500 147.0000 81.6000 ;
	    RECT 150.6000 81.4500 151.8000 81.6000 ;
	    RECT 145.8000 80.5500 151.8000 81.4500 ;
	    RECT 145.8000 80.4000 147.0000 80.5500 ;
	    RECT 150.6000 80.4000 151.8000 80.5500 ;
	    RECT 155.4000 80.4000 156.6000 81.6000 ;
	    RECT 162.3000 81.3000 162.6000 81.6000 ;
	    RECT 168.3000 81.3000 169.2000 84.3000 ;
	    RECT 174.6000 83.7000 175.8000 89.7000 ;
	    RECT 170.1000 82.2000 171.3000 83.4000 ;
	    RECT 172.2000 82.8000 175.8000 83.7000 ;
	    RECT 177.0000 83.7000 178.2000 89.7000 ;
	    RECT 179.4000 84.6000 180.9000 89.7000 ;
	    RECT 183.6000 84.3000 186.0000 89.7000 ;
	    RECT 188.7000 84.6000 190.2000 89.7000 ;
	    RECT 177.0000 82.8000 180.6000 83.7000 ;
	    RECT 172.2000 82.5000 173.4000 82.8000 ;
	    RECT 179.4000 82.5000 180.6000 82.8000 ;
	    RECT 162.3000 81.0000 163.5000 81.3000 ;
	    RECT 162.3000 80.4000 166.8000 81.0000 ;
	    RECT 162.6000 80.1000 166.8000 80.4000 ;
	    RECT 165.6000 79.8000 166.8000 80.1000 ;
	    RECT 167.7000 80.4000 169.2000 81.3000 ;
	    RECT 170.4000 81.6000 171.3000 82.2000 ;
	    RECT 181.5000 82.2000 182.7000 83.4000 ;
	    RECT 181.5000 81.6000 182.4000 82.2000 ;
	    RECT 170.4000 80.4000 171.6000 81.6000 ;
	    RECT 173.4000 80.4000 173.7000 81.6000 ;
	    RECT 177.0000 80.4000 178.2000 81.6000 ;
	    RECT 179.1000 80.4000 179.4000 81.6000 ;
	    RECT 181.2000 80.4000 182.4000 81.6000 ;
	    RECT 183.6000 81.3000 184.5000 84.3000 ;
	    RECT 191.4000 83.7000 192.6000 89.7000 ;
	    RECT 185.4000 82.2000 187.8000 83.4000 ;
	    RECT 188.7000 82.8000 192.6000 83.7000 ;
	    RECT 188.7000 82.5000 189.9000 82.8000 ;
	    RECT 190.2000 81.3000 190.5000 81.6000 ;
	    RECT 183.6000 80.4000 185.1000 81.3000 ;
	    RECT 189.3000 81.0000 190.5000 81.3000 ;
	    RECT 167.7000 79.5000 168.6000 80.4000 ;
	    RECT 184.2000 79.5000 185.1000 80.4000 ;
	    RECT 186.0000 80.4000 190.5000 81.0000 ;
	    RECT 191.4000 80.4000 192.6000 81.6000 ;
	    RECT 186.0000 80.1000 190.2000 80.4000 ;
	    RECT 186.0000 79.8000 187.2000 80.1000 ;
	    RECT 114.6000 77.4000 115.8000 78.6000 ;
	    RECT 114.6000 76.2000 115.8000 76.5000 ;
	    RECT 117.0000 75.3000 117.9000 79.5000 ;
	    RECT 124.2000 77.4000 125.4000 78.6000 ;
	    RECT 115.5000 74.1000 118.2000 75.3000 ;
	    RECT 115.5000 63.3000 116.7000 74.1000 ;
	    RECT 119.4000 63.3000 120.6000 75.3000 ;
	    RECT 121.8000 74.4000 123.0000 75.6000 ;
	    RECT 121.8000 73.2000 123.0000 73.5000 ;
	    RECT 121.8000 63.3000 123.0000 69.3000 ;
	    RECT 124.2000 63.3000 125.4000 76.5000 ;
	    RECT 126.6000 63.3000 127.8000 69.3000 ;
	    RECT 129.0000 63.3000 130.2000 69.3000 ;
	    RECT 131.4000 63.3000 132.6000 79.5000 ;
	    RECT 143.4000 77.4000 144.6000 78.6000 ;
	    RECT 148.2000 78.4500 149.4000 78.6000 ;
	    RECT 145.9500 77.5500 149.4000 78.4500 ;
	    RECT 141.0000 63.3000 142.2000 69.3000 ;
	    RECT 143.4000 63.3000 144.6000 76.5000 ;
	    RECT 145.9500 75.6000 146.8500 77.5500 ;
	    RECT 148.2000 77.4000 149.4000 77.5500 ;
	    RECT 148.2000 76.2000 149.4000 76.5000 ;
	    RECT 145.8000 74.4000 147.0000 75.6000 ;
	    RECT 150.6000 75.3000 151.5000 79.5000 ;
	    RECT 149.1000 74.1000 151.8000 75.3000 ;
	    RECT 145.8000 73.2000 147.0000 73.5000 ;
	    RECT 145.8000 63.3000 147.0000 69.3000 ;
	    RECT 149.1000 63.3000 150.3000 74.1000 ;
	    RECT 153.0000 63.3000 154.2000 75.3000 ;
	    RECT 155.4000 63.3000 156.6000 79.5000 ;
	    RECT 163.5000 78.3000 164.7000 78.6000 ;
	    RECT 163.5000 77.4000 165.9000 78.3000 ;
	    RECT 167.4000 77.4000 168.6000 78.6000 ;
	    RECT 184.2000 77.4000 185.4000 78.6000 ;
	    RECT 188.1000 78.3000 189.3000 78.6000 ;
	    RECT 186.9000 77.4000 189.3000 78.3000 ;
	    RECT 164.7000 77.1000 165.9000 77.4000 ;
	    RECT 186.9000 77.1000 188.1000 77.4000 ;
	    RECT 167.7000 75.3000 168.6000 76.5000 ;
	    RECT 184.2000 75.3000 185.1000 76.5000 ;
	    RECT 160.2000 74.4000 164.1000 75.3000 ;
	    RECT 157.8000 63.3000 159.0000 69.3000 ;
	    RECT 160.2000 63.3000 161.4000 74.4000 ;
	    RECT 162.9000 74.1000 164.1000 74.4000 ;
	    RECT 162.6000 63.3000 164.1000 73.2000 ;
	    RECT 166.8000 63.3000 169.2000 75.3000 ;
	    RECT 172.2000 74.4000 175.8000 75.3000 ;
	    RECT 172.2000 74.1000 173.4000 74.4000 ;
	    RECT 171.9000 63.3000 173.4000 73.2000 ;
	    RECT 174.6000 63.3000 175.8000 74.4000 ;
	    RECT 177.0000 74.4000 180.6000 75.3000 ;
	    RECT 177.0000 63.3000 178.2000 74.4000 ;
	    RECT 179.4000 74.1000 180.6000 74.4000 ;
	    RECT 179.4000 63.3000 180.9000 73.2000 ;
	    RECT 183.6000 63.3000 186.0000 75.3000 ;
	    RECT 188.7000 74.4000 192.6000 75.3000 ;
	    RECT 188.7000 74.1000 189.9000 74.4000 ;
	    RECT 188.7000 63.3000 190.2000 73.2000 ;
	    RECT 191.4000 63.3000 192.6000 74.4000 ;
	    RECT 0.6000 60.6000 193.8000 62.4000 ;
	    RECT 1.8000 48.6000 3.0000 59.7000 ;
	    RECT 4.2000 49.8000 5.7000 59.7000 ;
	    RECT 4.5000 48.6000 5.7000 48.9000 ;
	    RECT 1.8000 47.7000 5.7000 48.6000 ;
	    RECT 8.4000 47.7000 10.8000 59.7000 ;
	    RECT 13.5000 49.8000 15.0000 59.7000 ;
	    RECT 13.8000 48.6000 15.0000 48.9000 ;
	    RECT 16.2000 48.6000 17.4000 59.7000 ;
	    RECT 13.8000 47.7000 17.4000 48.6000 ;
	    RECT 18.6000 47.7000 19.8000 59.7000 ;
	    RECT 21.0000 49.5000 22.2000 59.7000 ;
	    RECT 23.4000 48.6000 24.6000 59.7000 ;
	    RECT 21.3000 47.7000 24.6000 48.6000 ;
	    RECT 25.8000 48.6000 27.0000 59.7000 ;
	    RECT 28.2000 49.8000 29.7000 59.7000 ;
	    RECT 28.5000 48.6000 29.7000 48.9000 ;
	    RECT 25.8000 47.7000 29.7000 48.6000 ;
	    RECT 32.4000 47.7000 34.8000 59.7000 ;
	    RECT 37.5000 49.8000 39.0000 59.7000 ;
	    RECT 37.8000 48.6000 39.0000 48.9000 ;
	    RECT 40.2000 48.6000 41.4000 59.7000 ;
	    RECT 42.6000 53.7000 43.8000 59.7000 ;
	    RECT 37.8000 47.7000 41.4000 48.6000 ;
	    RECT 9.3000 46.5000 10.2000 47.7000 ;
	    RECT 6.3000 45.6000 7.5000 45.9000 ;
	    RECT 5.1000 44.7000 7.5000 45.6000 ;
	    RECT 5.1000 44.4000 6.3000 44.7000 ;
	    RECT 9.0000 44.4000 10.2000 45.6000 ;
	    RECT 18.6000 44.4000 19.5000 47.7000 ;
	    RECT 21.3000 46.8000 22.2000 47.7000 ;
	    RECT 20.4000 45.6000 22.2000 46.8000 ;
	    RECT 33.3000 46.5000 34.2000 47.7000 ;
	    RECT 30.3000 45.6000 31.5000 45.9000 ;
	    RECT 18.6000 43.5000 19.8000 44.4000 ;
	    RECT 7.2000 42.9000 8.4000 43.2000 ;
	    RECT 4.2000 42.6000 8.4000 42.9000 ;
	    RECT 3.9000 42.0000 8.4000 42.6000 ;
	    RECT 9.3000 42.6000 10.2000 43.5000 ;
	    RECT 3.9000 41.7000 5.1000 42.0000 ;
	    RECT 9.3000 41.7000 10.8000 42.6000 ;
	    RECT 3.9000 41.4000 4.2000 41.7000 ;
	    RECT 4.5000 40.2000 5.7000 40.5000 ;
	    RECT 1.8000 39.3000 5.7000 40.2000 ;
	    RECT 6.6000 39.6000 9.0000 40.8000 ;
	    RECT 1.8000 33.3000 3.0000 39.3000 ;
	    RECT 9.9000 38.7000 10.8000 41.7000 ;
	    RECT 12.0000 41.4000 13.2000 42.6000 ;
	    RECT 15.0000 41.4000 15.3000 42.6000 ;
	    RECT 12.0000 40.8000 12.9000 41.4000 ;
	    RECT 11.7000 39.6000 12.9000 40.8000 ;
	    RECT 21.3000 41.1000 22.2000 45.6000 ;
	    RECT 23.4000 44.4000 24.6000 45.6000 ;
	    RECT 29.1000 44.7000 31.5000 45.6000 ;
	    RECT 29.1000 44.4000 30.3000 44.7000 ;
	    RECT 33.0000 44.4000 34.2000 45.6000 ;
	    RECT 45.0000 43.5000 46.2000 59.7000 ;
	    RECT 47.4000 53.7000 48.6000 59.7000 ;
	    RECT 49.8000 46.5000 51.0000 59.7000 ;
	    RECT 52.2000 53.7000 53.4000 59.7000 ;
	    RECT 61.8000 53.7000 63.0000 59.7000 ;
	    RECT 52.2000 49.5000 53.4000 49.8000 ;
	    RECT 61.8000 49.5000 63.0000 49.8000 ;
	    RECT 52.2000 47.4000 53.4000 48.6000 ;
	    RECT 61.8000 47.4000 63.0000 48.6000 ;
	    RECT 49.8000 44.4000 51.0000 45.6000 ;
	    RECT 52.3500 45.4500 53.2500 47.4000 ;
	    RECT 64.2000 46.5000 65.4000 59.7000 ;
	    RECT 66.6000 53.7000 67.8000 59.7000 ;
	    RECT 69.0000 53.7000 70.2000 59.7000 ;
	    RECT 69.0000 49.5000 70.2000 49.8000 ;
	    RECT 69.0000 47.4000 70.2000 48.6000 ;
	    RECT 71.4000 46.5000 72.6000 59.7000 ;
	    RECT 73.8000 53.7000 75.0000 59.7000 ;
	    RECT 76.2000 47.7000 77.4000 59.7000 ;
	    RECT 80.1000 48.9000 81.3000 59.7000 ;
	    RECT 78.6000 47.7000 81.3000 48.9000 ;
	    RECT 64.2000 45.4500 65.4000 45.6000 ;
	    RECT 52.3500 44.5500 65.4000 45.4500 ;
	    RECT 64.2000 44.4000 65.4000 44.5500 ;
	    RECT 71.4000 44.4000 72.6000 45.6000 ;
	    RECT 78.9000 43.5000 79.8000 47.7000 ;
	    RECT 81.0000 46.5000 82.2000 46.8000 ;
	    RECT 81.0000 44.4000 82.2000 45.6000 ;
	    RECT 83.4000 43.5000 84.6000 59.7000 ;
	    RECT 85.8000 53.7000 87.0000 59.7000 ;
	    RECT 88.2000 43.5000 89.4000 59.7000 ;
	    RECT 90.6000 53.7000 91.8000 59.7000 ;
	    RECT 93.0000 53.7000 94.2000 59.7000 ;
	    RECT 95.4000 46.5000 96.6000 59.7000 ;
	    RECT 97.8000 53.7000 99.0000 59.7000 ;
	    RECT 97.8000 49.5000 99.0000 49.8000 ;
	    RECT 97.8000 47.4000 99.0000 48.6000 ;
	    RECT 95.4000 44.4000 96.6000 45.6000 ;
	    RECT 100.2000 43.5000 101.4000 59.7000 ;
	    RECT 102.6000 53.7000 103.8000 59.7000 ;
	    RECT 105.0000 53.7000 106.2000 59.7000 ;
	    RECT 105.0000 49.5000 106.2000 49.8000 ;
	    RECT 105.0000 47.4000 106.2000 48.6000 ;
	    RECT 107.4000 46.5000 108.6000 59.7000 ;
	    RECT 109.8000 53.7000 111.0000 59.7000 ;
	    RECT 109.8000 50.4000 111.0000 51.6000 ;
	    RECT 102.6000 45.4500 103.8000 45.6000 ;
	    RECT 107.4000 45.4500 108.6000 45.6000 ;
	    RECT 102.6000 44.5500 108.6000 45.4500 ;
	    RECT 109.9500 45.4500 110.8500 50.4000 ;
	    RECT 112.2000 47.7000 113.4000 59.7000 ;
	    RECT 114.6000 48.3000 115.8000 59.7000 ;
	    RECT 117.0000 53.7000 118.2000 59.7000 ;
	    RECT 119.4000 53.7000 120.6000 59.7000 ;
	    RECT 121.8000 53.7000 123.0000 59.7000 ;
	    RECT 112.2000 46.5000 113.1000 47.7000 ;
	    RECT 117.0000 47.4000 117.9000 53.7000 ;
	    RECT 121.8000 47.4000 123.0000 48.6000 ;
	    RECT 114.3000 46.5000 117.9000 47.4000 ;
	    RECT 112.2000 45.4500 113.4000 45.6000 ;
	    RECT 109.9500 44.5500 113.4000 45.4500 ;
	    RECT 102.6000 44.4000 103.8000 44.5500 ;
	    RECT 107.4000 44.4000 108.6000 44.5500 ;
	    RECT 112.2000 44.4000 113.4000 44.5500 ;
	    RECT 23.4000 43.2000 24.6000 43.5000 ;
	    RECT 31.2000 42.9000 32.4000 43.2000 ;
	    RECT 28.2000 42.6000 32.4000 42.9000 ;
	    RECT 25.8000 41.4000 27.0000 42.6000 ;
	    RECT 27.9000 42.0000 32.4000 42.6000 ;
	    RECT 33.3000 42.6000 34.2000 43.5000 ;
	    RECT 27.9000 41.7000 29.1000 42.0000 ;
	    RECT 33.3000 41.7000 34.8000 42.6000 ;
	    RECT 27.9000 41.4000 28.2000 41.7000 ;
	    RECT 13.8000 40.2000 15.0000 40.5000 ;
	    RECT 13.8000 39.3000 17.4000 40.2000 ;
	    RECT 4.2000 33.3000 5.7000 38.4000 ;
	    RECT 8.4000 33.3000 10.8000 38.7000 ;
	    RECT 13.5000 33.3000 15.0000 38.4000 ;
	    RECT 16.2000 33.3000 17.4000 39.3000 ;
	    RECT 18.6000 33.3000 19.8000 40.5000 ;
	    RECT 21.3000 40.2000 24.6000 41.1000 ;
	    RECT 28.5000 40.2000 29.7000 40.5000 ;
	    RECT 21.0000 33.3000 22.2000 39.3000 ;
	    RECT 23.4000 33.3000 24.6000 40.2000 ;
	    RECT 25.8000 39.3000 29.7000 40.2000 ;
	    RECT 30.6000 39.6000 33.0000 40.8000 ;
	    RECT 25.8000 33.3000 27.0000 39.3000 ;
	    RECT 33.9000 38.7000 34.8000 41.7000 ;
	    RECT 36.0000 41.4000 37.2000 42.6000 ;
	    RECT 39.0000 41.4000 39.3000 42.6000 ;
	    RECT 40.2000 41.4000 41.4000 42.6000 ;
	    RECT 45.0000 42.4500 46.2000 42.6000 ;
	    RECT 47.4000 42.4500 48.6000 42.6000 ;
	    RECT 45.0000 41.5500 48.6000 42.4500 ;
	    RECT 45.0000 41.4000 46.2000 41.5500 ;
	    RECT 47.4000 41.4000 48.6000 41.5500 ;
	    RECT 36.0000 40.8000 36.9000 41.4000 ;
	    RECT 35.7000 39.6000 36.9000 40.8000 ;
	    RECT 37.8000 40.2000 39.0000 40.5000 ;
	    RECT 37.8000 39.3000 41.4000 40.2000 ;
	    RECT 28.2000 33.3000 29.7000 38.4000 ;
	    RECT 32.4000 33.3000 34.8000 38.7000 ;
	    RECT 37.5000 33.3000 39.0000 38.4000 ;
	    RECT 40.2000 33.3000 41.4000 39.3000 ;
	    RECT 42.6000 38.4000 43.8000 39.6000 ;
	    RECT 42.6000 37.2000 43.8000 37.5000 ;
	    RECT 42.6000 33.3000 43.8000 36.3000 ;
	    RECT 45.0000 33.3000 46.2000 40.5000 ;
	    RECT 47.4000 40.2000 48.6000 40.5000 ;
	    RECT 49.8000 39.3000 51.0000 43.5000 ;
	    RECT 64.2000 39.3000 65.4000 43.5000 ;
	    RECT 66.6000 41.4000 67.8000 42.6000 ;
	    RECT 66.6000 40.2000 67.8000 40.5000 ;
	    RECT 71.4000 39.3000 72.6000 43.5000 ;
	    RECT 73.8000 42.4500 75.0000 42.6000 ;
	    RECT 73.8000 41.5500 77.2500 42.4500 ;
	    RECT 73.8000 41.4000 75.0000 41.5500 ;
	    RECT 73.8000 40.2000 75.0000 40.5000 ;
	    RECT 76.3500 39.6000 77.2500 41.5500 ;
	    RECT 78.6000 41.4000 79.8000 42.6000 ;
	    RECT 81.0000 42.4500 82.2000 42.6000 ;
	    RECT 83.4000 42.4500 84.6000 42.6000 ;
	    RECT 81.0000 41.5500 84.6000 42.4500 ;
	    RECT 81.0000 41.4000 82.2000 41.5500 ;
	    RECT 83.4000 41.4000 84.6000 41.5500 ;
	    RECT 85.8000 42.4500 87.0000 42.6000 ;
	    RECT 88.2000 42.4500 89.4000 42.6000 ;
	    RECT 85.8000 41.5500 89.4000 42.4500 ;
	    RECT 85.8000 41.4000 87.0000 41.5500 ;
	    RECT 88.2000 41.4000 89.4000 41.5500 ;
	    RECT 93.0000 41.4000 94.2000 42.6000 ;
	    RECT 47.4000 33.3000 48.6000 39.3000 ;
	    RECT 49.8000 38.4000 52.5000 39.3000 ;
	    RECT 51.3000 33.3000 52.5000 38.4000 ;
	    RECT 62.7000 38.4000 65.4000 39.3000 ;
	    RECT 62.7000 33.3000 63.9000 38.4000 ;
	    RECT 66.6000 33.3000 67.8000 39.3000 ;
	    RECT 69.9000 38.4000 72.6000 39.3000 ;
	    RECT 69.9000 33.3000 71.1000 38.4000 ;
	    RECT 73.8000 33.3000 75.0000 39.3000 ;
	    RECT 76.2000 38.4000 77.4000 39.6000 ;
	    RECT 76.2000 37.2000 77.4000 37.5000 ;
	    RECT 78.9000 36.3000 79.8000 40.5000 ;
	    RECT 76.2000 33.3000 77.4000 36.3000 ;
	    RECT 78.6000 33.3000 79.8000 36.3000 ;
	    RECT 81.0000 33.3000 82.2000 36.3000 ;
	    RECT 83.4000 33.3000 84.6000 40.5000 ;
	    RECT 85.8000 37.2000 87.0000 37.5000 ;
	    RECT 85.8000 33.3000 87.0000 36.3000 ;
	    RECT 88.2000 33.3000 89.4000 40.5000 ;
	    RECT 93.0000 40.2000 94.2000 40.5000 ;
	    RECT 95.4000 39.3000 96.6000 43.5000 ;
	    RECT 97.8000 42.4500 99.0000 42.6000 ;
	    RECT 100.2000 42.4500 101.4000 42.6000 ;
	    RECT 97.8000 41.5500 101.4000 42.4500 ;
	    RECT 97.8000 41.4000 99.0000 41.5500 ;
	    RECT 100.2000 41.4000 101.4000 41.5500 ;
	    RECT 90.6000 37.2000 91.8000 37.5000 ;
	    RECT 90.6000 33.3000 91.8000 36.3000 ;
	    RECT 93.0000 33.3000 94.2000 39.3000 ;
	    RECT 95.4000 38.4000 98.1000 39.3000 ;
	    RECT 96.9000 33.3000 98.1000 38.4000 ;
	    RECT 100.2000 33.3000 101.4000 40.5000 ;
	    RECT 102.6000 38.4000 103.8000 39.6000 ;
	    RECT 107.4000 39.3000 108.6000 43.5000 ;
	    RECT 109.8000 41.4000 111.0000 42.6000 ;
	    RECT 109.8000 40.2000 111.0000 40.5000 ;
	    RECT 112.2000 39.3000 113.1000 43.5000 ;
	    RECT 114.3000 41.4000 115.2000 46.5000 ;
	    RECT 117.0000 44.4000 118.2000 45.6000 ;
	    RECT 121.9500 45.4500 122.8500 47.4000 ;
	    RECT 124.2000 46.5000 125.4000 59.7000 ;
	    RECT 126.6000 53.7000 127.8000 59.7000 ;
	    RECT 129.0000 53.7000 130.2000 59.7000 ;
	    RECT 126.6000 49.5000 127.8000 49.8000 ;
	    RECT 129.0000 49.5000 130.2000 49.8000 ;
	    RECT 126.6000 47.4000 127.8000 48.6000 ;
	    RECT 129.0000 47.4000 130.2000 48.6000 ;
	    RECT 124.2000 45.4500 125.4000 45.6000 ;
	    RECT 121.9500 44.5500 125.4000 45.4500 ;
	    RECT 126.7500 45.4500 127.6500 47.4000 ;
	    RECT 131.4000 46.5000 132.6000 59.7000 ;
	    RECT 133.8000 53.7000 135.0000 59.7000 ;
	    RECT 143.4000 53.7000 144.6000 59.7000 ;
	    RECT 143.4000 49.5000 144.6000 49.8000 ;
	    RECT 143.4000 47.4000 144.6000 48.6000 ;
	    RECT 145.8000 46.5000 147.0000 59.7000 ;
	    RECT 148.2000 53.7000 149.4000 59.7000 ;
	    RECT 150.6000 53.7000 151.8000 59.7000 ;
	    RECT 131.4000 45.4500 132.6000 45.6000 ;
	    RECT 126.7500 44.5500 132.6000 45.4500 ;
	    RECT 124.2000 44.4000 125.4000 44.5500 ;
	    RECT 131.4000 44.4000 132.6000 44.5500 ;
	    RECT 145.8000 45.4500 147.0000 45.6000 ;
	    RECT 150.6000 45.4500 151.8000 45.6000 ;
	    RECT 145.8000 44.5500 151.8000 45.4500 ;
	    RECT 145.8000 44.4000 147.0000 44.5500 ;
	    RECT 150.6000 44.4000 151.8000 44.5500 ;
	    RECT 119.4000 43.5000 120.6000 43.8000 ;
	    RECT 153.0000 43.5000 154.2000 59.7000 ;
	    RECT 155.4000 53.7000 156.6000 59.7000 ;
	    RECT 157.8000 46.5000 159.0000 59.7000 ;
	    RECT 160.2000 53.7000 161.4000 59.7000 ;
	    RECT 160.2000 49.5000 161.4000 49.8000 ;
	    RECT 160.2000 47.4000 161.4000 48.6000 ;
	    RECT 157.8000 44.4000 159.0000 45.6000 ;
	    RECT 162.6000 43.5000 163.8000 59.7000 ;
	    RECT 165.0000 53.7000 166.2000 59.7000 ;
	    RECT 167.4000 48.6000 168.6000 59.7000 ;
	    RECT 169.8000 49.8000 171.3000 59.7000 ;
	    RECT 169.8000 48.6000 171.0000 48.9000 ;
	    RECT 167.4000 47.7000 171.0000 48.6000 ;
	    RECT 174.0000 47.7000 176.4000 59.7000 ;
	    RECT 179.1000 49.8000 180.6000 59.7000 ;
	    RECT 179.1000 48.6000 180.3000 48.9000 ;
	    RECT 181.8000 48.6000 183.0000 59.7000 ;
	    RECT 179.1000 47.7000 183.0000 48.6000 ;
	    RECT 184.2000 48.6000 185.4000 59.7000 ;
	    RECT 186.6000 49.5000 187.8000 59.7000 ;
	    RECT 184.2000 47.7000 187.5000 48.6000 ;
	    RECT 189.0000 47.7000 190.2000 59.7000 ;
	    RECT 174.6000 46.5000 175.5000 47.7000 ;
	    RECT 186.6000 46.8000 187.5000 47.7000 ;
	    RECT 177.3000 45.6000 178.5000 45.9000 ;
	    RECT 186.6000 45.6000 188.4000 46.8000 ;
	    RECT 172.2000 45.4500 173.4000 45.6000 ;
	    RECT 174.6000 45.4500 175.8000 45.6000 ;
	    RECT 172.2000 44.5500 175.8000 45.4500 ;
	    RECT 177.3000 44.7000 179.7000 45.6000 ;
	    RECT 172.2000 44.4000 173.4000 44.5500 ;
	    RECT 174.6000 44.4000 175.8000 44.5500 ;
	    RECT 178.5000 44.4000 179.7000 44.7000 ;
	    RECT 184.2000 44.4000 185.4000 45.6000 ;
	    RECT 117.0000 43.2000 117.9000 43.5000 ;
	    RECT 116.4000 42.3000 117.9000 43.2000 ;
	    RECT 116.4000 42.0000 117.6000 42.3000 ;
	    RECT 119.4000 41.4000 120.6000 42.6000 ;
	    RECT 121.8000 41.4000 123.0000 42.6000 ;
	    RECT 114.0000 41.1000 115.2000 41.4000 ;
	    RECT 114.0000 40.5000 118.5000 41.1000 ;
	    RECT 114.0000 40.2000 120.3000 40.5000 ;
	    RECT 121.8000 40.2000 123.0000 40.5000 ;
	    RECT 117.6000 39.6000 120.3000 40.2000 ;
	    RECT 119.4000 39.3000 120.3000 39.6000 ;
	    RECT 124.2000 39.3000 125.4000 43.5000 ;
	    RECT 131.4000 39.3000 132.6000 43.5000 ;
	    RECT 133.8000 42.4500 135.0000 42.6000 ;
	    RECT 143.4000 42.4500 144.6000 42.6000 ;
	    RECT 133.8000 41.5500 144.6000 42.4500 ;
	    RECT 133.8000 41.4000 135.0000 41.5500 ;
	    RECT 143.4000 41.4000 144.6000 41.5500 ;
	    RECT 133.8000 40.2000 135.0000 40.5000 ;
	    RECT 145.8000 39.3000 147.0000 43.5000 ;
	    RECT 148.2000 41.4000 149.4000 42.6000 ;
	    RECT 153.0000 42.4500 154.2000 42.6000 ;
	    RECT 155.4000 42.4500 156.6000 42.6000 ;
	    RECT 153.0000 41.5500 156.6000 42.4500 ;
	    RECT 153.0000 41.4000 154.2000 41.5500 ;
	    RECT 155.4000 41.4000 156.6000 41.5500 ;
	    RECT 148.2000 40.2000 149.4000 40.5000 ;
	    RECT 105.9000 38.4000 108.6000 39.3000 ;
	    RECT 102.6000 37.2000 103.8000 37.5000 ;
	    RECT 102.6000 33.3000 103.8000 36.3000 ;
	    RECT 105.9000 33.3000 107.1000 38.4000 ;
	    RECT 109.8000 33.3000 111.0000 39.3000 ;
	    RECT 112.2000 37.8000 114.3000 39.3000 ;
	    RECT 113.1000 33.3000 114.3000 37.8000 ;
	    RECT 115.5000 33.3000 116.7000 39.0000 ;
	    RECT 119.4000 33.3000 120.6000 39.3000 ;
	    RECT 121.8000 33.3000 123.0000 39.3000 ;
	    RECT 124.2000 38.4000 126.9000 39.3000 ;
	    RECT 125.7000 33.3000 126.9000 38.4000 ;
	    RECT 129.9000 38.4000 132.6000 39.3000 ;
	    RECT 129.9000 33.3000 131.1000 38.4000 ;
	    RECT 133.8000 33.3000 135.0000 39.3000 ;
	    RECT 144.3000 38.4000 147.0000 39.3000 ;
	    RECT 144.3000 33.3000 145.5000 38.4000 ;
	    RECT 148.2000 33.3000 149.4000 39.3000 ;
	    RECT 150.6000 38.4000 151.8000 39.6000 ;
	    RECT 150.6000 37.2000 151.8000 37.5000 ;
	    RECT 150.6000 33.3000 151.8000 36.3000 ;
	    RECT 153.0000 33.3000 154.2000 40.5000 ;
	    RECT 155.4000 40.2000 156.6000 40.5000 ;
	    RECT 157.8000 39.3000 159.0000 43.5000 ;
	    RECT 174.6000 42.6000 175.5000 43.5000 ;
	    RECT 184.2000 43.2000 185.4000 43.5000 ;
	    RECT 162.6000 41.4000 163.8000 42.6000 ;
	    RECT 167.4000 41.4000 168.6000 42.6000 ;
	    RECT 169.5000 41.4000 169.8000 42.6000 ;
	    RECT 171.6000 41.4000 172.8000 42.6000 ;
	    RECT 171.9000 40.8000 172.8000 41.4000 ;
	    RECT 174.0000 41.7000 175.5000 42.6000 ;
	    RECT 176.4000 42.9000 177.6000 43.2000 ;
	    RECT 176.4000 42.6000 180.6000 42.9000 ;
	    RECT 176.4000 42.0000 180.9000 42.6000 ;
	    RECT 179.7000 41.7000 180.9000 42.0000 ;
	    RECT 155.4000 33.3000 156.6000 39.3000 ;
	    RECT 157.8000 38.4000 160.5000 39.3000 ;
	    RECT 159.3000 33.3000 160.5000 38.4000 ;
	    RECT 162.6000 33.3000 163.8000 40.5000 ;
	    RECT 169.8000 40.2000 171.0000 40.5000 ;
	    RECT 167.4000 39.3000 171.0000 40.2000 ;
	    RECT 171.9000 39.6000 173.1000 40.8000 ;
	    RECT 165.0000 37.2000 166.2000 37.5000 ;
	    RECT 165.0000 33.3000 166.2000 36.3000 ;
	    RECT 167.4000 33.3000 168.6000 39.3000 ;
	    RECT 174.0000 38.7000 174.9000 41.7000 ;
	    RECT 180.6000 41.4000 180.9000 41.7000 ;
	    RECT 181.8000 41.4000 183.0000 42.6000 ;
	    RECT 186.6000 41.1000 187.5000 45.6000 ;
	    RECT 189.3000 44.4000 190.2000 47.7000 ;
	    RECT 189.0000 43.5000 190.2000 44.4000 ;
	    RECT 175.8000 39.6000 178.2000 40.8000 ;
	    RECT 179.1000 40.2000 180.3000 40.5000 ;
	    RECT 184.2000 40.2000 187.5000 41.1000 ;
	    RECT 179.1000 39.3000 183.0000 40.2000 ;
	    RECT 169.8000 33.3000 171.3000 38.4000 ;
	    RECT 174.0000 33.3000 176.4000 38.7000 ;
	    RECT 179.1000 33.3000 180.6000 38.4000 ;
	    RECT 181.8000 33.3000 183.0000 39.3000 ;
	    RECT 184.2000 33.3000 185.4000 40.2000 ;
	    RECT 186.6000 33.3000 187.8000 39.3000 ;
	    RECT 189.0000 33.3000 190.2000 40.5000 ;
	    RECT 0.6000 30.6000 193.8000 32.4000 ;
	    RECT 1.8000 26.7000 3.0000 29.7000 ;
	    RECT 1.8000 25.5000 3.0000 25.8000 ;
	    RECT 4.2000 22.5000 5.4000 29.7000 ;
	    RECT 6.6000 26.7000 7.8000 29.7000 ;
	    RECT 6.6000 25.5000 7.8000 25.8000 ;
	    RECT 9.0000 22.5000 10.2000 29.7000 ;
	    RECT 11.4000 26.7000 12.6000 29.7000 ;
	    RECT 13.8000 26.7000 15.0000 29.7000 ;
	    RECT 16.2000 26.7000 17.4000 29.7000 ;
	    RECT 13.8000 22.5000 14.7000 26.7000 ;
	    RECT 16.2000 25.5000 17.4000 25.8000 ;
	    RECT 16.2000 23.4000 17.4000 24.6000 ;
	    RECT 18.6000 23.7000 19.8000 29.7000 ;
	    RECT 22.5000 24.6000 23.7000 29.7000 ;
	    RECT 25.8000 26.7000 27.0000 29.7000 ;
	    RECT 25.8000 25.5000 27.0000 25.8000 ;
	    RECT 21.0000 23.7000 23.7000 24.6000 ;
	    RECT 4.2000 20.4000 5.4000 21.6000 ;
	    RECT 9.0000 21.4500 10.2000 21.6000 ;
	    RECT 9.0000 20.5500 12.4500 21.4500 ;
	    RECT 9.0000 20.4000 10.2000 20.5500 ;
	    RECT 1.8000 3.3000 3.0000 9.3000 ;
	    RECT 4.2000 3.3000 5.4000 19.5000 ;
	    RECT 6.6000 3.3000 7.8000 9.3000 ;
	    RECT 9.0000 3.3000 10.2000 19.5000 ;
	    RECT 11.5500 18.6000 12.4500 20.5500 ;
	    RECT 13.8000 20.4000 15.0000 21.6000 ;
	    RECT 16.3500 21.4500 17.2500 23.4000 ;
	    RECT 18.6000 22.5000 19.8000 22.8000 ;
	    RECT 18.6000 21.4500 19.8000 21.6000 ;
	    RECT 16.3500 20.5500 19.8000 21.4500 ;
	    RECT 18.6000 20.4000 19.8000 20.5500 ;
	    RECT 21.0000 19.5000 22.2000 23.7000 ;
	    RECT 25.8000 23.4000 27.0000 24.6000 ;
	    RECT 28.2000 22.5000 29.4000 29.7000 ;
	    RECT 30.6000 23.7000 31.8000 29.7000 ;
	    RECT 34.5000 24.6000 35.7000 29.7000 ;
	    RECT 33.0000 23.7000 35.7000 24.6000 ;
	    RECT 38.7000 24.6000 39.9000 29.7000 ;
	    RECT 38.7000 23.7000 41.4000 24.6000 ;
	    RECT 42.6000 23.7000 43.8000 29.7000 ;
	    RECT 45.0000 26.7000 46.2000 29.7000 ;
	    RECT 45.0000 25.5000 46.2000 25.8000 ;
	    RECT 30.6000 22.5000 31.8000 22.8000 ;
	    RECT 28.2000 21.4500 29.4000 21.6000 ;
	    RECT 30.6000 21.4500 31.8000 21.6000 ;
	    RECT 28.2000 20.5500 31.8000 21.4500 ;
	    RECT 28.2000 20.4000 29.4000 20.5500 ;
	    RECT 30.6000 20.4000 31.8000 20.5500 ;
	    RECT 33.0000 19.5000 34.2000 23.7000 ;
	    RECT 40.2000 19.5000 41.4000 23.7000 ;
	    RECT 45.0000 23.4000 46.2000 24.6000 ;
	    RECT 42.6000 22.5000 43.8000 22.8000 ;
	    RECT 47.4000 22.5000 48.6000 29.7000 ;
	    RECT 57.0000 23.7000 58.2000 29.7000 ;
	    RECT 60.9000 24.0000 62.1000 29.7000 ;
	    RECT 63.3000 25.2000 64.5000 29.7000 ;
	    RECT 63.3000 23.7000 65.4000 25.2000 ;
	    RECT 67.5000 24.6000 68.7000 29.7000 ;
	    RECT 67.5000 23.7000 70.2000 24.6000 ;
	    RECT 71.4000 23.7000 72.6000 29.7000 ;
	    RECT 74.7000 24.6000 75.9000 29.7000 ;
	    RECT 74.7000 23.7000 77.4000 24.6000 ;
	    RECT 78.6000 23.7000 79.8000 29.7000 ;
	    RECT 57.3000 23.4000 58.2000 23.7000 ;
	    RECT 57.3000 22.8000 60.0000 23.4000 ;
	    RECT 57.3000 22.5000 63.6000 22.8000 ;
	    RECT 59.1000 21.9000 63.6000 22.5000 ;
	    RECT 62.4000 21.6000 63.6000 21.9000 ;
	    RECT 42.6000 20.4000 43.8000 21.6000 ;
	    RECT 47.4000 21.4500 48.6000 21.6000 ;
	    RECT 54.6000 21.4500 55.8000 21.6000 ;
	    RECT 47.4000 20.5500 55.8000 21.4500 ;
	    RECT 47.4000 20.4000 48.6000 20.5500 ;
	    RECT 54.6000 20.4000 55.8000 20.5500 ;
	    RECT 57.0000 20.4000 58.2000 21.6000 ;
	    RECT 60.0000 20.7000 61.2000 21.0000 ;
	    RECT 59.7000 19.8000 61.2000 20.7000 ;
	    RECT 59.7000 19.5000 60.6000 19.8000 ;
	    RECT 11.4000 17.4000 12.6000 18.6000 ;
	    RECT 11.4000 16.2000 12.6000 16.5000 ;
	    RECT 13.8000 15.3000 14.7000 19.5000 ;
	    RECT 21.0000 17.4000 22.2000 18.6000 ;
	    RECT 12.3000 14.1000 15.0000 15.3000 ;
	    RECT 12.3000 3.3000 13.5000 14.1000 ;
	    RECT 16.2000 3.3000 17.4000 15.3000 ;
	    RECT 18.6000 3.3000 19.8000 9.3000 ;
	    RECT 21.0000 3.3000 22.2000 16.5000 ;
	    RECT 23.4000 14.4000 24.6000 15.6000 ;
	    RECT 23.4000 13.2000 24.6000 13.5000 ;
	    RECT 23.4000 3.3000 24.6000 9.3000 ;
	    RECT 25.8000 3.3000 27.0000 9.3000 ;
	    RECT 28.2000 3.3000 29.4000 19.5000 ;
	    RECT 33.0000 17.4000 34.2000 18.6000 ;
	    RECT 40.2000 18.4500 41.4000 18.6000 ;
	    RECT 35.5500 17.5500 41.4000 18.4500 ;
	    RECT 30.6000 3.3000 31.8000 9.3000 ;
	    RECT 33.0000 3.3000 34.2000 16.5000 ;
	    RECT 35.5500 15.6000 36.4500 17.5500 ;
	    RECT 40.2000 17.4000 41.4000 17.5500 ;
	    RECT 35.4000 14.4000 36.6000 15.6000 ;
	    RECT 37.8000 14.4000 39.0000 15.6000 ;
	    RECT 35.4000 13.2000 36.6000 13.5000 ;
	    RECT 37.8000 13.2000 39.0000 13.5000 ;
	    RECT 35.4000 3.3000 36.6000 9.3000 ;
	    RECT 37.8000 3.3000 39.0000 9.3000 ;
	    RECT 40.2000 3.3000 41.4000 16.5000 ;
	    RECT 42.6000 3.3000 43.8000 9.3000 ;
	    RECT 45.0000 3.3000 46.2000 9.3000 ;
	    RECT 47.4000 3.3000 48.6000 19.5000 ;
	    RECT 57.0000 19.2000 58.2000 19.5000 ;
	    RECT 59.4000 17.4000 60.6000 18.6000 ;
	    RECT 62.4000 16.5000 63.3000 21.6000 ;
	    RECT 64.5000 19.5000 65.4000 23.7000 ;
	    RECT 69.0000 19.5000 70.2000 23.7000 ;
	    RECT 71.4000 22.5000 72.6000 22.8000 ;
	    RECT 71.4000 20.4000 72.6000 21.6000 ;
	    RECT 76.2000 19.5000 77.4000 23.7000 ;
	    RECT 81.0000 22.8000 82.2000 29.7000 ;
	    RECT 83.4000 23.7000 84.6000 29.7000 ;
	    RECT 78.6000 22.5000 79.8000 22.8000 ;
	    RECT 81.0000 21.9000 84.3000 22.8000 ;
	    RECT 85.8000 22.5000 87.0000 29.7000 ;
	    RECT 88.2000 22.5000 89.4000 29.7000 ;
	    RECT 90.6000 23.7000 91.8000 29.7000 ;
	    RECT 93.0000 22.8000 94.2000 29.7000 ;
	    RECT 95.4000 23.7000 96.6000 29.7000 ;
	    RECT 97.8000 24.6000 99.3000 29.7000 ;
	    RECT 102.0000 24.3000 104.4000 29.7000 ;
	    RECT 107.1000 24.6000 108.6000 29.7000 ;
	    RECT 95.4000 22.8000 99.0000 23.7000 ;
	    RECT 78.6000 20.4000 79.8000 21.6000 ;
	    RECT 81.0000 19.5000 82.2000 19.8000 ;
	    RECT 64.2000 18.4500 65.4000 18.6000 ;
	    RECT 69.0000 18.4500 70.2000 18.6000 ;
	    RECT 76.2000 18.4500 77.4000 18.6000 ;
	    RECT 81.0000 18.4500 82.2000 18.6000 ;
	    RECT 64.2000 17.5500 67.6500 18.4500 ;
	    RECT 64.2000 17.4000 65.4000 17.5500 ;
	    RECT 59.7000 15.6000 63.3000 16.5000 ;
	    RECT 59.7000 9.3000 60.6000 15.6000 ;
	    RECT 64.5000 15.3000 65.4000 16.5000 ;
	    RECT 66.7500 15.6000 67.6500 17.5500 ;
	    RECT 69.0000 17.5500 74.8500 18.4500 ;
	    RECT 69.0000 17.4000 70.2000 17.5500 ;
	    RECT 57.0000 3.3000 58.2000 9.3000 ;
	    RECT 59.4000 3.3000 60.6000 9.3000 ;
	    RECT 61.8000 3.3000 63.0000 14.7000 ;
	    RECT 64.2000 3.3000 65.4000 15.3000 ;
	    RECT 66.6000 14.4000 67.8000 15.6000 ;
	    RECT 66.6000 13.2000 67.8000 13.5000 ;
	    RECT 66.6000 3.3000 67.8000 9.3000 ;
	    RECT 69.0000 3.3000 70.2000 16.5000 ;
	    RECT 73.9500 15.6000 74.8500 17.5500 ;
	    RECT 76.2000 17.5500 82.2000 18.4500 ;
	    RECT 76.2000 17.4000 77.4000 17.5500 ;
	    RECT 81.0000 17.4000 82.2000 17.5500 ;
	    RECT 83.4000 17.4000 84.3000 21.9000 ;
	    RECT 90.9000 21.9000 94.2000 22.8000 ;
	    RECT 97.8000 22.5000 99.0000 22.8000 ;
	    RECT 99.9000 22.2000 101.1000 23.4000 ;
	    RECT 85.8000 18.6000 87.0000 19.5000 ;
	    RECT 73.8000 14.4000 75.0000 15.6000 ;
	    RECT 73.8000 13.2000 75.0000 13.5000 ;
	    RECT 71.4000 3.3000 72.6000 9.3000 ;
	    RECT 73.8000 3.3000 75.0000 9.3000 ;
	    RECT 76.2000 3.3000 77.4000 16.5000 ;
	    RECT 83.4000 16.2000 85.2000 17.4000 ;
	    RECT 83.4000 15.3000 84.3000 16.2000 ;
	    RECT 86.1000 15.3000 87.0000 18.6000 ;
	    RECT 81.0000 14.4000 84.3000 15.3000 ;
	    RECT 78.6000 3.3000 79.8000 9.3000 ;
	    RECT 81.0000 3.3000 82.2000 14.4000 ;
	    RECT 83.4000 3.3000 84.6000 13.5000 ;
	    RECT 85.8000 3.3000 87.0000 15.3000 ;
	    RECT 88.2000 18.6000 89.4000 19.5000 ;
	    RECT 88.2000 15.3000 89.1000 18.6000 ;
	    RECT 90.9000 17.4000 91.8000 21.9000 ;
	    RECT 99.9000 21.6000 100.8000 22.2000 ;
	    RECT 95.4000 20.4000 96.6000 21.6000 ;
	    RECT 97.5000 20.4000 97.8000 21.6000 ;
	    RECT 99.6000 20.4000 100.8000 21.6000 ;
	    RECT 102.0000 21.3000 102.9000 24.3000 ;
	    RECT 109.8000 23.7000 111.0000 29.7000 ;
	    RECT 103.8000 22.2000 106.2000 23.4000 ;
	    RECT 107.1000 22.8000 111.0000 23.7000 ;
	    RECT 112.2000 23.7000 113.4000 29.7000 ;
	    RECT 114.6000 24.6000 116.1000 29.7000 ;
	    RECT 118.8000 24.3000 121.2000 29.7000 ;
	    RECT 123.9000 24.6000 125.4000 29.7000 ;
	    RECT 112.2000 22.8000 116.1000 23.7000 ;
	    RECT 107.1000 22.5000 108.3000 22.8000 ;
	    RECT 114.9000 22.5000 116.1000 22.8000 ;
	    RECT 117.0000 22.2000 119.4000 23.4000 ;
	    RECT 108.6000 21.3000 108.9000 21.6000 ;
	    RECT 102.0000 20.4000 103.5000 21.3000 ;
	    RECT 107.7000 21.0000 108.9000 21.3000 ;
	    RECT 93.0000 19.5000 94.2000 19.8000 ;
	    RECT 102.6000 19.5000 103.5000 20.4000 ;
	    RECT 104.4000 20.4000 108.9000 21.0000 ;
	    RECT 109.8000 20.4000 111.0000 21.6000 ;
	    RECT 114.3000 21.3000 114.6000 21.6000 ;
	    RECT 120.3000 21.3000 121.2000 24.3000 ;
	    RECT 126.6000 23.7000 127.8000 29.7000 ;
	    RECT 122.1000 22.2000 123.3000 23.4000 ;
	    RECT 124.2000 22.8000 127.8000 23.7000 ;
	    RECT 124.2000 22.5000 125.4000 22.8000 ;
	    RECT 129.0000 22.5000 130.2000 29.7000 ;
	    RECT 131.4000 26.7000 132.6000 29.7000 ;
	    RECT 131.4000 25.5000 132.6000 25.8000 ;
	    RECT 131.4000 24.4500 132.6000 24.6000 ;
	    RECT 138.6000 24.4500 139.8000 24.6000 ;
	    RECT 131.4000 23.5500 139.8000 24.4500 ;
	    RECT 141.0000 23.7000 142.2000 29.7000 ;
	    RECT 144.9000 24.6000 146.1000 29.7000 ;
	    RECT 148.2000 26.7000 149.4000 29.7000 ;
	    RECT 150.6000 26.7000 151.8000 29.7000 ;
	    RECT 153.0000 26.7000 154.2000 29.7000 ;
	    RECT 143.4000 23.7000 146.1000 24.6000 ;
	    RECT 131.4000 23.4000 132.6000 23.5500 ;
	    RECT 138.6000 23.4000 139.8000 23.5500 ;
	    RECT 141.0000 22.5000 142.2000 22.8000 ;
	    RECT 114.3000 21.0000 115.5000 21.3000 ;
	    RECT 114.3000 20.4000 118.8000 21.0000 ;
	    RECT 104.4000 20.1000 108.6000 20.4000 ;
	    RECT 114.6000 20.1000 118.8000 20.4000 ;
	    RECT 104.4000 19.8000 105.6000 20.1000 ;
	    RECT 117.6000 19.8000 118.8000 20.1000 ;
	    RECT 119.7000 20.4000 121.2000 21.3000 ;
	    RECT 122.4000 21.6000 123.3000 22.2000 ;
	    RECT 122.4000 20.4000 123.6000 21.6000 ;
	    RECT 125.4000 20.4000 125.7000 21.6000 ;
	    RECT 129.0000 20.4000 130.2000 21.6000 ;
	    RECT 141.0000 20.4000 142.2000 21.6000 ;
	    RECT 119.7000 19.5000 120.6000 20.4000 ;
	    RECT 143.4000 19.5000 144.6000 23.7000 ;
	    RECT 150.6000 22.5000 151.5000 26.7000 ;
	    RECT 153.0000 25.5000 154.2000 25.8000 ;
	    RECT 153.0000 23.4000 154.2000 24.6000 ;
	    RECT 155.4000 22.5000 156.6000 29.7000 ;
	    RECT 157.8000 26.7000 159.0000 29.7000 ;
	    RECT 157.8000 25.5000 159.0000 25.8000 ;
	    RECT 160.2000 22.5000 161.4000 29.7000 ;
	    RECT 162.6000 26.7000 163.8000 29.7000 ;
	    RECT 162.6000 25.5000 163.8000 25.8000 ;
	    RECT 165.0000 23.7000 166.2000 29.7000 ;
	    RECT 167.4000 24.6000 168.9000 29.7000 ;
	    RECT 171.6000 24.3000 174.0000 29.7000 ;
	    RECT 176.7000 24.6000 178.2000 29.7000 ;
	    RECT 165.0000 22.8000 168.9000 23.7000 ;
	    RECT 167.7000 22.5000 168.9000 22.8000 ;
	    RECT 169.8000 22.2000 172.2000 23.4000 ;
	    RECT 145.8000 21.4500 147.0000 21.6000 ;
	    RECT 150.6000 21.4500 151.8000 21.6000 ;
	    RECT 145.8000 20.5500 151.8000 21.4500 ;
	    RECT 145.8000 20.4000 147.0000 20.5500 ;
	    RECT 150.6000 20.4000 151.8000 20.5500 ;
	    RECT 153.0000 21.4500 154.2000 21.6000 ;
	    RECT 155.4000 21.4500 156.6000 21.6000 ;
	    RECT 153.0000 20.5500 156.6000 21.4500 ;
	    RECT 153.0000 20.4000 154.2000 20.5500 ;
	    RECT 155.4000 20.4000 156.6000 20.5500 ;
	    RECT 160.2000 20.4000 161.4000 21.6000 ;
	    RECT 167.1000 21.3000 167.4000 21.6000 ;
	    RECT 173.1000 21.3000 174.0000 24.3000 ;
	    RECT 179.4000 23.7000 180.6000 29.7000 ;
	    RECT 174.9000 22.2000 176.1000 23.4000 ;
	    RECT 177.0000 22.8000 180.6000 23.7000 ;
	    RECT 181.8000 22.8000 183.0000 29.7000 ;
	    RECT 184.2000 23.7000 185.4000 29.7000 ;
	    RECT 177.0000 22.5000 178.2000 22.8000 ;
	    RECT 167.1000 21.0000 168.3000 21.3000 ;
	    RECT 167.1000 20.4000 171.6000 21.0000 ;
	    RECT 167.4000 20.1000 171.6000 20.4000 ;
	    RECT 170.4000 19.8000 171.6000 20.1000 ;
	    RECT 172.5000 20.4000 174.0000 21.3000 ;
	    RECT 175.2000 21.6000 176.1000 22.2000 ;
	    RECT 181.8000 21.9000 185.1000 22.8000 ;
	    RECT 186.6000 22.5000 187.8000 29.7000 ;
	    RECT 175.2000 20.4000 176.4000 21.6000 ;
	    RECT 178.2000 20.4000 178.5000 21.6000 ;
	    RECT 172.5000 19.5000 173.4000 20.4000 ;
	    RECT 181.8000 19.5000 183.0000 19.8000 ;
	    RECT 93.0000 18.4500 94.2000 18.6000 ;
	    RECT 102.6000 18.4500 103.8000 18.6000 ;
	    RECT 93.0000 17.5500 103.8000 18.4500 ;
	    RECT 106.5000 18.3000 107.7000 18.6000 ;
	    RECT 93.0000 17.4000 94.2000 17.5500 ;
	    RECT 102.6000 17.4000 103.8000 17.5500 ;
	    RECT 105.3000 17.4000 107.7000 18.3000 ;
	    RECT 115.5000 18.3000 116.7000 18.6000 ;
	    RECT 115.5000 17.4000 117.9000 18.3000 ;
	    RECT 119.4000 17.4000 120.6000 18.6000 ;
	    RECT 90.0000 16.2000 91.8000 17.4000 ;
	    RECT 105.3000 17.1000 106.5000 17.4000 ;
	    RECT 116.7000 17.1000 117.9000 17.4000 ;
	    RECT 90.9000 15.3000 91.8000 16.2000 ;
	    RECT 102.6000 15.3000 103.5000 16.5000 ;
	    RECT 119.7000 15.3000 120.6000 16.5000 ;
	    RECT 88.2000 3.3000 89.4000 15.3000 ;
	    RECT 90.9000 14.4000 94.2000 15.3000 ;
	    RECT 90.6000 3.3000 91.8000 13.5000 ;
	    RECT 93.0000 3.3000 94.2000 14.4000 ;
	    RECT 95.4000 14.4000 99.0000 15.3000 ;
	    RECT 95.4000 3.3000 96.6000 14.4000 ;
	    RECT 97.8000 14.1000 99.0000 14.4000 ;
	    RECT 97.8000 3.3000 99.3000 13.2000 ;
	    RECT 102.0000 3.3000 104.4000 15.3000 ;
	    RECT 107.1000 14.4000 111.0000 15.3000 ;
	    RECT 107.1000 14.1000 108.3000 14.4000 ;
	    RECT 107.1000 3.3000 108.6000 13.2000 ;
	    RECT 109.8000 3.3000 111.0000 14.4000 ;
	    RECT 112.2000 14.4000 116.1000 15.3000 ;
	    RECT 112.2000 3.3000 113.4000 14.4000 ;
	    RECT 114.9000 14.1000 116.1000 14.4000 ;
	    RECT 114.6000 3.3000 116.1000 13.2000 ;
	    RECT 118.8000 3.3000 121.2000 15.3000 ;
	    RECT 124.2000 14.4000 127.8000 15.3000 ;
	    RECT 124.2000 14.1000 125.4000 14.4000 ;
	    RECT 123.9000 3.3000 125.4000 13.2000 ;
	    RECT 126.6000 3.3000 127.8000 14.4000 ;
	    RECT 129.0000 3.3000 130.2000 19.5000 ;
	    RECT 131.4000 18.4500 132.6000 18.6000 ;
	    RECT 143.4000 18.4500 144.6000 18.6000 ;
	    RECT 148.2000 18.4500 149.4000 18.6000 ;
	    RECT 131.4000 17.5500 144.6000 18.4500 ;
	    RECT 131.4000 17.4000 132.6000 17.5500 ;
	    RECT 143.4000 17.4000 144.6000 17.5500 ;
	    RECT 145.9500 17.5500 149.4000 18.4500 ;
	    RECT 131.4000 3.3000 132.6000 9.3000 ;
	    RECT 141.0000 3.3000 142.2000 9.3000 ;
	    RECT 143.4000 3.3000 144.6000 16.5000 ;
	    RECT 145.9500 15.6000 146.8500 17.5500 ;
	    RECT 148.2000 17.4000 149.4000 17.5500 ;
	    RECT 148.2000 16.2000 149.4000 16.5000 ;
	    RECT 145.8000 14.4000 147.0000 15.6000 ;
	    RECT 150.6000 15.3000 151.5000 19.5000 ;
	    RECT 149.1000 14.1000 151.8000 15.3000 ;
	    RECT 145.8000 13.2000 147.0000 13.5000 ;
	    RECT 145.8000 3.3000 147.0000 9.3000 ;
	    RECT 149.1000 3.3000 150.3000 14.1000 ;
	    RECT 153.0000 3.3000 154.2000 15.3000 ;
	    RECT 155.4000 3.3000 156.6000 19.5000 ;
	    RECT 157.8000 3.3000 159.0000 9.3000 ;
	    RECT 160.2000 3.3000 161.4000 19.5000 ;
	    RECT 168.3000 18.3000 169.5000 18.6000 ;
	    RECT 172.2000 18.4500 173.4000 18.6000 ;
	    RECT 174.6000 18.4500 175.8000 18.6000 ;
	    RECT 168.3000 17.4000 170.7000 18.3000 ;
	    RECT 172.2000 17.5500 175.8000 18.4500 ;
	    RECT 172.2000 17.4000 173.4000 17.5500 ;
	    RECT 174.6000 17.4000 175.8000 17.5500 ;
	    RECT 181.8000 17.4000 183.0000 18.6000 ;
	    RECT 184.2000 17.4000 185.1000 21.9000 ;
	    RECT 186.6000 18.6000 187.8000 19.5000 ;
	    RECT 169.5000 17.1000 170.7000 17.4000 ;
	    RECT 172.5000 15.3000 173.4000 16.5000 ;
	    RECT 184.2000 16.2000 186.0000 17.4000 ;
	    RECT 184.2000 15.3000 185.1000 16.2000 ;
	    RECT 186.9000 15.3000 187.8000 18.6000 ;
	    RECT 165.0000 14.4000 168.9000 15.3000 ;
	    RECT 162.6000 3.3000 163.8000 9.3000 ;
	    RECT 165.0000 3.3000 166.2000 14.4000 ;
	    RECT 167.7000 14.1000 168.9000 14.4000 ;
	    RECT 167.4000 3.3000 168.9000 13.2000 ;
	    RECT 171.6000 3.3000 174.0000 15.3000 ;
	    RECT 177.0000 14.4000 180.6000 15.3000 ;
	    RECT 177.0000 14.1000 178.2000 14.4000 ;
	    RECT 176.7000 3.3000 178.2000 13.2000 ;
	    RECT 179.4000 3.3000 180.6000 14.4000 ;
	    RECT 181.8000 14.4000 185.1000 15.3000 ;
	    RECT 181.8000 3.3000 183.0000 14.4000 ;
	    RECT 184.2000 3.3000 185.4000 13.5000 ;
	    RECT 186.6000 3.3000 187.8000 15.3000 ;
	    RECT 0.6000 0.6000 193.8000 2.4000 ;
         LAYER metal2 ;
	    RECT 133.2000 90.6000 140.4000 92.4000 ;
	    RECT 11.7000 83.4000 12.9000 83.7000 ;
	    RECT 11.7000 82.5000 20.1000 83.4000 ;
	    RECT 21.0000 82.5000 22.2000 83.7000 ;
	    RECT 9.0000 77.4000 10.2000 78.6000 ;
	    RECT 11.7000 75.3000 12.6000 82.5000 ;
	    RECT 13.8000 82.2000 15.0000 82.5000 ;
	    RECT 18.9000 82.2000 20.1000 82.5000 ;
	    RECT 21.3000 81.3000 22.2000 82.5000 ;
	    RECT 59.4000 82.5000 60.6000 83.7000 ;
	    RECT 68.7000 83.4000 69.9000 83.7000 ;
	    RECT 61.5000 82.5000 69.9000 83.4000 ;
	    RECT 13.8000 80.4000 22.2000 81.3000 ;
	    RECT 33.0000 80.4000 34.2000 81.6000 ;
	    RECT 49.8000 80.4000 51.0000 81.6000 ;
	    RECT 59.4000 81.3000 60.3000 82.5000 ;
	    RECT 61.5000 82.2000 62.7000 82.5000 ;
	    RECT 66.6000 82.2000 67.8000 82.5000 ;
	    RECT 59.4000 80.4000 67.8000 81.3000 ;
	    RECT 13.8000 78.3000 14.7000 80.4000 ;
	    RECT 13.5000 77.1000 14.7000 78.3000 ;
	    RECT 16.2000 77.4000 17.4000 78.6000 ;
	    RECT 21.3000 75.3000 22.2000 80.4000 ;
	    RECT 33.1500 78.6000 34.0500 80.4000 ;
	    RECT 49.9500 78.6000 50.8500 80.4000 ;
	    RECT 33.0000 77.4000 34.2000 78.6000 ;
	    RECT 49.8000 77.4000 51.0000 78.6000 ;
	    RECT 11.7000 74.1000 12.9000 75.3000 ;
	    RECT 21.0000 74.1000 22.2000 75.3000 ;
	    RECT 59.4000 75.3000 60.3000 80.4000 ;
	    RECT 66.9000 78.3000 67.8000 80.4000 ;
	    RECT 66.9000 77.1000 68.1000 78.3000 ;
	    RECT 69.0000 75.3000 69.9000 82.5000 ;
	    RECT 76.5000 83.4000 77.7000 83.7000 ;
	    RECT 76.5000 82.5000 84.9000 83.4000 ;
	    RECT 85.8000 82.5000 87.0000 83.7000 ;
	    RECT 102.6000 83.4000 103.8000 84.6000 ;
	    RECT 119.4000 83.4000 120.6000 84.6000 ;
	    RECT 124.2000 83.4000 125.4000 84.6000 ;
	    RECT 129.0000 83.4000 130.2000 84.6000 ;
	    RECT 153.0000 83.4000 154.2000 84.6000 ;
	    RECT 162.9000 83.4000 164.1000 83.7000 ;
	    RECT 71.4000 80.4000 72.6000 81.6000 ;
	    RECT 59.4000 74.1000 60.6000 75.3000 ;
	    RECT 68.7000 74.1000 69.9000 75.3000 ;
	    RECT 71.5500 72.6000 72.4500 80.4000 ;
	    RECT 76.5000 75.3000 77.4000 82.5000 ;
	    RECT 78.6000 82.2000 79.8000 82.5000 ;
	    RECT 83.7000 82.2000 84.9000 82.5000 ;
	    RECT 86.1000 81.3000 87.0000 82.5000 ;
	    RECT 102.7500 81.6000 103.6500 83.4000 ;
	    RECT 78.6000 80.4000 87.0000 81.3000 ;
	    RECT 90.6000 80.4000 91.8000 81.6000 ;
	    RECT 102.6000 80.4000 103.8000 81.6000 ;
	    RECT 107.4000 80.4000 108.6000 81.6000 ;
	    RECT 121.8000 81.4500 123.0000 81.6000 ;
	    RECT 124.3500 81.4500 125.2500 83.4000 ;
	    RECT 121.8000 80.5500 125.2500 81.4500 ;
	    RECT 121.8000 80.4000 123.0000 80.5500 ;
	    RECT 141.0000 80.4000 142.2000 81.6000 ;
	    RECT 145.8000 80.4000 147.0000 81.6000 ;
	    RECT 78.6000 78.3000 79.5000 80.4000 ;
	    RECT 78.3000 77.1000 79.5000 78.3000 ;
	    RECT 81.0000 77.4000 82.2000 78.6000 ;
	    RECT 76.5000 74.1000 77.7000 75.3000 ;
	    RECT 81.1500 72.6000 82.0500 77.4000 ;
	    RECT 86.1000 75.3000 87.0000 80.4000 ;
	    RECT 90.7500 78.6000 91.6500 80.4000 ;
	    RECT 90.6000 77.4000 91.8000 78.6000 ;
	    RECT 95.4000 77.4000 96.6000 78.6000 ;
	    RECT 97.8000 77.4000 99.0000 78.6000 ;
	    RECT 105.0000 77.4000 106.2000 78.6000 ;
	    RECT 85.8000 74.1000 87.0000 75.3000 ;
	    RECT 95.5500 72.6000 96.4500 77.4000 ;
	    RECT 97.9500 75.6000 98.8500 77.4000 ;
	    RECT 107.5500 75.6000 108.4500 80.4000 ;
	    RECT 124.2000 77.4000 125.4000 78.6000 ;
	    RECT 97.8000 74.4000 99.0000 75.6000 ;
	    RECT 107.4000 74.4000 108.6000 75.6000 ;
	    RECT 121.8000 74.4000 123.0000 75.6000 ;
	    RECT 121.9500 72.6000 122.8500 74.4000 ;
	    RECT 71.4000 71.4000 72.6000 72.6000 ;
	    RECT 81.0000 71.4000 82.2000 72.6000 ;
	    RECT 95.4000 71.4000 96.6000 72.6000 ;
	    RECT 121.8000 71.4000 123.0000 72.6000 ;
	    RECT 51.6000 60.6000 58.8000 62.4000 ;
	    RECT 105.0000 53.4000 106.2000 54.6000 ;
	    RECT 109.8000 53.4000 111.0000 54.6000 ;
	    RECT 4.5000 47.7000 5.7000 48.9000 ;
	    RECT 13.8000 47.7000 15.0000 48.9000 ;
	    RECT 4.5000 40.5000 5.4000 47.7000 ;
	    RECT 6.3000 44.7000 7.5000 45.9000 ;
	    RECT 6.6000 42.6000 7.5000 44.7000 ;
	    RECT 9.0000 44.4000 10.2000 45.6000 ;
	    RECT 14.1000 42.6000 15.0000 47.7000 ;
	    RECT 23.4000 47.4000 24.6000 48.6000 ;
	    RECT 28.5000 47.7000 29.7000 48.9000 ;
	    RECT 23.5500 45.6000 24.4500 47.4000 ;
	    RECT 23.4000 44.4000 24.6000 45.6000 ;
	    RECT 6.6000 41.7000 15.0000 42.6000 ;
	    RECT 6.6000 40.5000 7.8000 40.8000 ;
	    RECT 11.7000 40.5000 12.9000 40.8000 ;
	    RECT 14.1000 40.5000 15.0000 41.7000 ;
	    RECT 25.8000 41.4000 27.0000 42.6000 ;
	    RECT 4.5000 39.6000 12.9000 40.5000 ;
	    RECT 4.5000 39.3000 5.7000 39.6000 ;
	    RECT 13.8000 39.3000 15.0000 40.5000 ;
	    RECT 28.5000 40.5000 29.4000 47.7000 ;
	    RECT 33.0000 47.4000 34.2000 48.6000 ;
	    RECT 37.8000 47.7000 39.0000 48.9000 ;
	    RECT 105.1500 48.6000 106.0500 53.4000 ;
	    RECT 109.9500 51.6000 110.8500 53.4000 ;
	    RECT 109.8000 50.4000 111.0000 51.6000 ;
	    RECT 112.3500 50.5500 122.8500 51.4500 ;
	    RECT 30.3000 44.7000 31.5000 45.9000 ;
	    RECT 33.1500 45.6000 34.0500 47.4000 ;
	    RECT 30.6000 42.6000 31.5000 44.7000 ;
	    RECT 33.0000 44.4000 34.2000 45.6000 ;
	    RECT 38.1000 42.6000 39.0000 47.7000 ;
	    RECT 40.2000 47.4000 41.4000 48.6000 ;
	    RECT 49.8000 47.4000 51.0000 48.6000 ;
	    RECT 61.8000 48.4500 63.0000 48.6000 ;
	    RECT 59.5500 47.5500 63.0000 48.4500 ;
	    RECT 40.3500 42.6000 41.2500 47.4000 ;
	    RECT 49.9500 45.6000 50.8500 47.4000 ;
	    RECT 49.8000 44.4000 51.0000 45.6000 ;
	    RECT 30.6000 41.7000 39.0000 42.6000 ;
	    RECT 30.6000 40.5000 31.8000 40.8000 ;
	    RECT 35.7000 40.5000 36.9000 40.8000 ;
	    RECT 38.1000 40.5000 39.0000 41.7000 ;
	    RECT 40.2000 41.4000 41.4000 42.6000 ;
	    RECT 42.6000 41.4000 43.8000 42.6000 ;
	    RECT 28.5000 39.6000 36.9000 40.5000 ;
	    RECT 28.5000 39.3000 29.7000 39.6000 ;
	    RECT 37.8000 39.3000 39.0000 40.5000 ;
	    RECT 42.7500 39.6000 43.6500 41.4000 ;
	    RECT 42.6000 38.4000 43.8000 39.6000 ;
	    RECT 13.9500 26.5500 22.0500 27.4500 ;
	    RECT 4.2000 23.4000 5.4000 24.6000 ;
	    RECT 4.3500 21.6000 5.2500 23.4000 ;
	    RECT 13.9500 21.6000 14.8500 26.5500 ;
	    RECT 21.1500 24.6000 22.0500 26.5500 ;
	    RECT 16.2000 23.4000 17.4000 24.6000 ;
	    RECT 21.0000 23.4000 22.2000 24.6000 ;
	    RECT 25.8000 23.4000 27.0000 24.6000 ;
	    RECT 33.0000 23.4000 34.2000 24.6000 ;
	    RECT 4.2000 20.4000 5.4000 21.6000 ;
	    RECT 13.8000 20.4000 15.0000 21.6000 ;
	    RECT 33.1500 18.6000 34.0500 23.4000 ;
	    RECT 42.7500 21.6000 43.6500 38.4000 ;
	    RECT 45.0000 23.4000 46.2000 24.6000 ;
	    RECT 54.6000 23.4000 55.8000 24.6000 ;
	    RECT 54.7500 21.6000 55.6500 23.4000 ;
	    RECT 42.6000 20.4000 43.8000 21.6000 ;
	    RECT 54.6000 20.4000 55.8000 21.6000 ;
	    RECT 57.0000 20.4000 58.2000 21.6000 ;
	    RECT 57.1500 18.6000 58.0500 20.4000 ;
	    RECT 59.5500 18.6000 60.4500 47.5500 ;
	    RECT 61.8000 47.4000 63.0000 47.5500 ;
	    RECT 69.0000 47.4000 70.2000 48.6000 ;
	    RECT 71.4000 47.4000 72.6000 48.6000 ;
	    RECT 76.2000 47.4000 77.4000 48.6000 ;
	    RECT 81.0000 47.4000 82.2000 48.6000 ;
	    RECT 85.8000 47.4000 87.0000 48.6000 ;
	    RECT 97.8000 47.4000 99.0000 48.6000 ;
	    RECT 102.6000 47.4000 103.8000 48.6000 ;
	    RECT 105.0000 47.4000 106.2000 48.6000 ;
	    RECT 109.8000 47.4000 111.0000 48.6000 ;
	    RECT 66.6000 41.4000 67.8000 42.6000 ;
	    RECT 69.1500 42.4500 70.0500 47.4000 ;
	    RECT 71.5500 45.6000 72.4500 47.4000 ;
	    RECT 71.4000 44.4000 72.6000 45.6000 ;
	    RECT 76.3500 45.4500 77.2500 47.4000 ;
	    RECT 81.1500 45.6000 82.0500 47.4000 ;
	    RECT 73.9500 44.5500 77.2500 45.4500 ;
	    RECT 73.9500 42.4500 74.8500 44.5500 ;
	    RECT 81.0000 44.4000 82.2000 45.6000 ;
	    RECT 85.9500 42.6000 86.8500 47.4000 ;
	    RECT 102.7500 45.6000 103.6500 47.4000 ;
	    RECT 95.4000 44.4000 96.6000 45.6000 ;
	    RECT 102.6000 44.4000 103.8000 45.6000 ;
	    RECT 69.1500 41.5500 74.8500 42.4500 ;
	    RECT 78.6000 41.4000 79.8000 42.6000 ;
	    RECT 81.0000 41.4000 82.2000 42.6000 ;
	    RECT 85.8000 41.4000 87.0000 42.6000 ;
	    RECT 93.0000 41.4000 94.2000 42.6000 ;
	    RECT 66.7500 30.6000 67.6500 41.4000 ;
	    RECT 76.2000 38.4000 77.4000 39.6000 ;
	    RECT 76.3500 36.6000 77.2500 38.4000 ;
	    RECT 81.1500 36.6000 82.0500 41.4000 ;
	    RECT 76.2000 35.4000 77.4000 36.6000 ;
	    RECT 81.0000 35.4000 82.2000 36.6000 ;
	    RECT 95.5500 30.6000 96.4500 44.4000 ;
	    RECT 109.9500 42.6000 110.8500 47.4000 ;
	    RECT 112.3500 42.6000 113.2500 50.5500 ;
	    RECT 121.9500 48.6000 122.8500 50.5500 ;
	    RECT 124.3500 48.6000 125.2500 77.4000 ;
	    RECT 141.1500 66.6000 142.0500 80.4000 ;
	    RECT 143.4000 77.4000 144.6000 78.6000 ;
	    RECT 141.0000 65.4000 142.2000 66.6000 ;
	    RECT 143.5500 60.6000 144.4500 77.4000 ;
	    RECT 126.6000 59.4000 127.8000 60.6000 ;
	    RECT 143.4000 59.4000 144.6000 60.6000 ;
	    RECT 114.7500 47.5500 120.4500 48.4500 ;
	    RECT 97.8000 41.4000 99.0000 42.6000 ;
	    RECT 102.6000 41.4000 103.8000 42.6000 ;
	    RECT 109.8000 41.4000 111.0000 42.6000 ;
	    RECT 112.2000 41.4000 113.4000 42.6000 ;
	    RECT 102.7500 39.6000 103.6500 41.4000 ;
	    RECT 102.6000 38.4000 103.8000 39.6000 ;
	    RECT 114.7500 36.6000 115.6500 47.5500 ;
	    RECT 117.0000 44.4000 118.2000 45.6000 ;
	    RECT 119.5500 45.4500 120.4500 47.5500 ;
	    RECT 121.8000 47.4000 123.0000 48.6000 ;
	    RECT 124.2000 47.4000 125.4000 48.6000 ;
	    RECT 126.7500 45.4500 127.6500 59.4000 ;
	    RECT 143.5500 48.6000 144.4500 59.4000 ;
	    RECT 129.0000 47.4000 130.2000 48.6000 ;
	    RECT 143.4000 47.4000 144.6000 48.6000 ;
	    RECT 119.5500 44.5500 122.8500 45.4500 ;
	    RECT 117.1500 39.4500 118.0500 44.4000 ;
	    RECT 121.9500 42.6000 122.8500 44.5500 ;
	    RECT 124.3500 44.5500 127.6500 45.4500 ;
	    RECT 119.4000 41.4000 120.6000 42.6000 ;
	    RECT 121.8000 41.4000 123.0000 42.6000 ;
	    RECT 124.3500 39.4500 125.2500 44.5500 ;
	    RECT 129.1500 42.6000 130.0500 47.4000 ;
	    RECT 129.0000 41.4000 130.2000 42.6000 ;
	    RECT 143.4000 42.4500 144.6000 42.6000 ;
	    RECT 145.9500 42.4500 146.8500 80.4000 ;
	    RECT 148.2000 77.4000 149.4000 78.6000 ;
	    RECT 148.3500 72.6000 149.2500 77.4000 ;
	    RECT 148.2000 71.4000 149.4000 72.6000 ;
	    RECT 153.1500 66.6000 154.0500 83.4000 ;
	    RECT 162.9000 82.5000 171.3000 83.4000 ;
	    RECT 172.2000 82.5000 173.4000 83.7000 ;
	    RECT 155.4000 80.4000 156.6000 81.6000 ;
	    RECT 155.5500 72.6000 156.4500 80.4000 ;
	    RECT 162.9000 75.3000 163.8000 82.5000 ;
	    RECT 165.0000 82.2000 166.2000 82.5000 ;
	    RECT 170.1000 82.2000 171.3000 82.5000 ;
	    RECT 172.5000 81.3000 173.4000 82.5000 ;
	    RECT 179.4000 82.5000 180.6000 83.7000 ;
	    RECT 188.7000 83.4000 189.9000 83.7000 ;
	    RECT 181.5000 82.5000 189.9000 83.4000 ;
	    RECT 165.0000 80.4000 173.4000 81.3000 ;
	    RECT 177.0000 80.4000 178.2000 81.6000 ;
	    RECT 179.4000 81.3000 180.3000 82.5000 ;
	    RECT 181.5000 82.2000 182.7000 82.5000 ;
	    RECT 186.6000 82.2000 187.8000 82.5000 ;
	    RECT 179.4000 80.4000 187.8000 81.3000 ;
	    RECT 165.0000 78.3000 165.9000 80.4000 ;
	    RECT 164.7000 77.1000 165.9000 78.3000 ;
	    RECT 167.4000 77.4000 168.6000 78.6000 ;
	    RECT 172.5000 75.3000 173.4000 80.4000 ;
	    RECT 162.9000 74.1000 164.1000 75.3000 ;
	    RECT 172.2000 74.1000 173.4000 75.3000 ;
	    RECT 155.4000 71.4000 156.6000 72.6000 ;
	    RECT 153.0000 65.4000 154.2000 66.6000 ;
	    RECT 162.6000 65.4000 163.8000 66.6000 ;
	    RECT 150.6000 53.4000 151.8000 54.6000 ;
	    RECT 160.2000 53.4000 161.4000 54.6000 ;
	    RECT 148.2000 47.4000 149.4000 48.6000 ;
	    RECT 148.3500 42.6000 149.2500 47.4000 ;
	    RECT 150.7500 45.6000 151.6500 53.4000 ;
	    RECT 160.3500 48.6000 161.2500 53.4000 ;
	    RECT 160.2000 47.4000 161.4000 48.6000 ;
	    RECT 150.6000 44.4000 151.8000 45.6000 ;
	    RECT 157.8000 44.4000 159.0000 45.6000 ;
	    RECT 143.4000 41.5500 146.8500 42.4500 ;
	    RECT 143.4000 41.4000 144.6000 41.5500 ;
	    RECT 148.2000 41.4000 149.4000 42.6000 ;
	    RECT 150.6000 41.4000 151.8000 42.6000 ;
	    RECT 117.1500 38.5500 125.2500 39.4500 ;
	    RECT 114.6000 35.4000 115.8000 36.6000 ;
	    RECT 126.6000 35.4000 127.8000 36.6000 ;
	    RECT 66.6000 29.4000 67.8000 30.6000 ;
	    RECT 71.4000 29.4000 72.6000 30.6000 ;
	    RECT 95.4000 29.4000 96.6000 30.6000 ;
	    RECT 71.5500 21.6000 72.4500 29.4000 ;
	    RECT 78.6000 23.4000 79.8000 24.6000 ;
	    RECT 78.7500 21.6000 79.6500 23.4000 ;
	    RECT 95.5500 21.6000 96.4500 29.4000 ;
	    RECT 97.8000 22.5000 99.0000 23.7000 ;
	    RECT 107.1000 23.4000 108.3000 23.7000 ;
	    RECT 99.9000 22.5000 108.3000 23.4000 ;
	    RECT 71.4000 20.4000 72.6000 21.6000 ;
	    RECT 78.6000 20.4000 79.8000 21.6000 ;
	    RECT 95.4000 20.4000 96.6000 21.6000 ;
	    RECT 97.8000 21.3000 98.7000 22.5000 ;
	    RECT 99.9000 22.2000 101.1000 22.5000 ;
	    RECT 105.0000 22.2000 106.2000 22.5000 ;
	    RECT 97.8000 20.4000 106.2000 21.3000 ;
	    RECT 11.4000 17.4000 12.6000 18.6000 ;
	    RECT 16.2000 17.4000 17.4000 18.6000 ;
	    RECT 21.0000 17.4000 22.2000 18.6000 ;
	    RECT 33.0000 17.4000 34.2000 18.6000 ;
	    RECT 37.8000 17.4000 39.0000 18.6000 ;
	    RECT 57.0000 17.4000 58.2000 18.6000 ;
	    RECT 59.4000 17.4000 60.6000 18.6000 ;
	    RECT 16.3500 15.4500 17.2500 17.4000 ;
	    RECT 37.9500 15.6000 38.8500 17.4000 ;
	    RECT 23.4000 15.4500 24.6000 15.6000 ;
	    RECT 16.3500 14.5500 24.6000 15.4500 ;
	    RECT 23.4000 14.4000 24.6000 14.5500 ;
	    RECT 37.8000 14.4000 39.0000 15.6000 ;
	    RECT 97.8000 15.3000 98.7000 20.4000 ;
	    RECT 105.3000 18.3000 106.2000 20.4000 ;
	    RECT 105.3000 17.1000 106.5000 18.3000 ;
	    RECT 107.4000 15.3000 108.3000 22.5000 ;
	    RECT 114.9000 23.4000 116.1000 23.7000 ;
	    RECT 114.9000 22.5000 123.3000 23.4000 ;
	    RECT 124.2000 22.5000 125.4000 23.7000 ;
	    RECT 109.8000 20.4000 111.0000 21.6000 ;
	    RECT 97.8000 14.1000 99.0000 15.3000 ;
	    RECT 107.1000 14.1000 108.3000 15.3000 ;
	    RECT 109.9500 12.4500 110.8500 20.4000 ;
	    RECT 114.9000 15.3000 115.8000 22.5000 ;
	    RECT 117.0000 22.2000 118.2000 22.5000 ;
	    RECT 122.1000 22.2000 123.3000 22.5000 ;
	    RECT 124.5000 21.3000 125.4000 22.5000 ;
	    RECT 117.0000 20.4000 125.4000 21.3000 ;
	    RECT 126.7500 21.4500 127.6500 35.4000 ;
	    RECT 129.1500 24.4500 130.0500 41.4000 ;
	    RECT 150.7500 39.6000 151.6500 41.4000 ;
	    RECT 150.6000 38.4000 151.8000 39.6000 ;
	    RECT 157.9500 36.6000 158.8500 44.4000 ;
	    RECT 162.7500 42.6000 163.6500 65.4000 ;
	    RECT 169.8000 47.7000 171.0000 48.9000 ;
	    RECT 177.1500 48.6000 178.0500 80.4000 ;
	    RECT 179.4000 75.3000 180.3000 80.4000 ;
	    RECT 184.2000 77.4000 185.4000 78.6000 ;
	    RECT 186.9000 78.3000 187.8000 80.4000 ;
	    RECT 179.4000 74.1000 180.6000 75.3000 ;
	    RECT 169.8000 42.6000 170.7000 47.7000 ;
	    RECT 177.0000 47.4000 178.2000 48.6000 ;
	    RECT 179.1000 47.7000 180.3000 48.9000 ;
	    RECT 172.2000 44.4000 173.4000 45.6000 ;
	    RECT 177.3000 44.7000 178.5000 45.9000 ;
	    RECT 177.3000 42.6000 178.2000 44.7000 ;
	    RECT 162.6000 41.4000 163.8000 42.6000 ;
	    RECT 167.4000 41.4000 168.6000 42.6000 ;
	    RECT 169.8000 41.7000 178.2000 42.6000 ;
	    RECT 167.5500 36.6000 168.4500 41.4000 ;
	    RECT 169.8000 40.5000 170.7000 41.7000 ;
	    RECT 171.9000 40.5000 173.1000 40.8000 ;
	    RECT 177.0000 40.5000 178.2000 40.8000 ;
	    RECT 179.4000 40.5000 180.3000 47.7000 ;
	    RECT 184.3500 48.4500 185.2500 77.4000 ;
	    RECT 186.9000 77.1000 188.1000 78.3000 ;
	    RECT 189.0000 75.3000 189.9000 82.5000 ;
	    RECT 191.4000 80.4000 192.6000 81.6000 ;
	    RECT 191.5500 78.6000 192.4500 80.4000 ;
	    RECT 191.4000 77.4000 192.6000 78.6000 ;
	    RECT 188.7000 74.1000 189.9000 75.3000 ;
	    RECT 184.3500 47.5500 187.6500 48.4500 ;
	    RECT 184.2000 44.4000 185.4000 45.6000 ;
	    RECT 184.3500 42.6000 185.2500 44.4000 ;
	    RECT 181.8000 41.4000 183.0000 42.6000 ;
	    RECT 184.2000 41.4000 185.4000 42.6000 ;
	    RECT 169.8000 39.3000 171.0000 40.5000 ;
	    RECT 171.9000 39.6000 180.3000 40.5000 ;
	    RECT 179.1000 39.3000 180.3000 39.6000 ;
	    RECT 157.8000 35.4000 159.0000 36.6000 ;
	    RECT 167.4000 35.4000 168.6000 36.6000 ;
	    RECT 181.9500 33.4500 182.8500 41.4000 ;
	    RECT 181.9500 32.5500 185.2500 33.4500 ;
	    RECT 133.2000 30.6000 140.4000 32.4000 ;
	    RECT 181.8000 29.4000 183.0000 30.6000 ;
	    RECT 129.1500 23.5500 132.4500 24.4500 ;
	    RECT 129.0000 21.4500 130.2000 21.6000 ;
	    RECT 126.7500 20.5500 130.2000 21.4500 ;
	    RECT 129.0000 20.4000 130.2000 20.5500 ;
	    RECT 117.0000 18.3000 117.9000 20.4000 ;
	    RECT 116.7000 17.1000 117.9000 18.3000 ;
	    RECT 119.4000 17.4000 120.6000 18.6000 ;
	    RECT 119.5500 15.4500 120.4500 17.4000 ;
	    RECT 114.9000 14.1000 116.1000 15.3000 ;
	    RECT 117.1500 14.5500 120.4500 15.4500 ;
	    RECT 124.5000 15.3000 125.4000 20.4000 ;
	    RECT 131.5500 18.6000 132.4500 23.5500 ;
	    RECT 138.6000 23.4000 139.8000 24.6000 ;
	    RECT 141.0000 23.4000 142.2000 24.6000 ;
	    RECT 153.0000 23.4000 154.2000 24.6000 ;
	    RECT 160.2000 23.4000 161.4000 24.6000 ;
	    RECT 167.7000 23.4000 168.9000 23.7000 ;
	    RECT 138.7500 18.6000 139.6500 23.4000 ;
	    RECT 141.1500 21.6000 142.0500 23.4000 ;
	    RECT 160.3500 21.6000 161.2500 23.4000 ;
	    RECT 167.7000 22.5000 176.1000 23.4000 ;
	    RECT 177.0000 22.5000 178.2000 23.7000 ;
	    RECT 141.0000 20.4000 142.2000 21.6000 ;
	    RECT 145.8000 21.4500 147.0000 21.6000 ;
	    RECT 143.5500 20.5500 147.0000 21.4500 ;
	    RECT 143.5500 18.6000 144.4500 20.5500 ;
	    RECT 145.8000 20.4000 147.0000 20.5500 ;
	    RECT 153.0000 20.4000 154.2000 21.6000 ;
	    RECT 160.2000 20.4000 161.4000 21.6000 ;
	    RECT 153.1500 18.6000 154.0500 20.4000 ;
	    RECT 131.4000 17.4000 132.6000 18.6000 ;
	    RECT 138.6000 17.4000 139.8000 18.6000 ;
	    RECT 143.4000 17.4000 144.6000 18.6000 ;
	    RECT 148.2000 17.4000 149.4000 18.6000 ;
	    RECT 153.0000 17.4000 154.2000 18.6000 ;
	    RECT 117.1500 12.4500 118.0500 14.5500 ;
	    RECT 124.2000 14.1000 125.4000 15.3000 ;
	    RECT 167.7000 15.3000 168.6000 22.5000 ;
	    RECT 169.8000 22.2000 171.0000 22.5000 ;
	    RECT 174.9000 22.2000 176.1000 22.5000 ;
	    RECT 177.3000 21.3000 178.2000 22.5000 ;
	    RECT 169.8000 20.4000 178.2000 21.3000 ;
	    RECT 169.8000 18.3000 170.7000 20.4000 ;
	    RECT 169.5000 17.1000 170.7000 18.3000 ;
	    RECT 174.6000 17.4000 175.8000 18.6000 ;
	    RECT 167.7000 14.1000 168.9000 15.3000 ;
	    RECT 174.7500 12.6000 175.6500 17.4000 ;
	    RECT 177.3000 15.3000 178.2000 20.4000 ;
	    RECT 181.9500 18.6000 182.8500 29.4000 ;
	    RECT 181.8000 17.4000 183.0000 18.6000 ;
	    RECT 184.3500 15.4500 185.2500 32.5500 ;
	    RECT 186.7500 30.6000 187.6500 47.5500 ;
	    RECT 186.6000 29.4000 187.8000 30.6000 ;
	    RECT 177.0000 14.1000 178.2000 15.3000 ;
	    RECT 179.5500 14.5500 185.2500 15.4500 ;
	    RECT 179.5500 12.6000 180.4500 14.5500 ;
	    RECT 109.9500 11.5500 118.0500 12.4500 ;
	    RECT 174.6000 11.4000 175.8000 12.6000 ;
	    RECT 179.4000 11.4000 180.6000 12.6000 ;
	    RECT 51.6000 0.6000 58.8000 2.4000 ;
         LAYER metal3 ;
	    RECT 133.2000 90.6000 140.4000 92.4000 ;
	    RECT 102.3000 84.7500 104.1000 84.9000 ;
	    RECT 119.1000 84.7500 120.9000 84.9000 ;
	    RECT 102.3000 83.2500 120.9000 84.7500 ;
	    RECT 102.3000 83.1000 104.1000 83.2500 ;
	    RECT 119.1000 83.1000 120.9000 83.2500 ;
	    RECT 123.9000 84.7500 125.7000 84.9000 ;
	    RECT 128.7000 84.7500 130.5000 84.9000 ;
	    RECT 123.9000 83.2500 130.5000 84.7500 ;
	    RECT 123.9000 83.1000 125.7000 83.2500 ;
	    RECT 128.7000 83.1000 130.5000 83.2500 ;
	    RECT 8.7000 78.7500 10.5000 78.9000 ;
	    RECT 15.9000 78.7500 17.7000 78.9000 ;
	    RECT 8.7000 77.2500 17.7000 78.7500 ;
	    RECT 8.7000 77.1000 10.5000 77.2500 ;
	    RECT 15.9000 77.1000 17.7000 77.2500 ;
	    RECT 32.7000 78.7500 34.5000 78.9000 ;
	    RECT 49.5000 78.7500 51.3000 78.9000 ;
	    RECT 90.3000 78.7500 92.1000 78.9000 ;
	    RECT 32.7000 77.2500 92.1000 78.7500 ;
	    RECT 32.7000 77.1000 34.5000 77.2500 ;
	    RECT 49.5000 77.1000 51.3000 77.2500 ;
	    RECT 90.3000 77.1000 92.1000 77.2500 ;
	    RECT 97.5000 78.7500 99.3000 78.9000 ;
	    RECT 104.7000 78.7500 106.5000 78.9000 ;
	    RECT 97.5000 77.2500 106.5000 78.7500 ;
	    RECT 97.5000 77.1000 99.3000 77.2500 ;
	    RECT 104.7000 77.1000 106.5000 77.2500 ;
	    RECT 167.1000 78.7500 168.9000 78.9000 ;
	    RECT 191.1000 78.7500 192.9000 78.9000 ;
	    RECT 167.1000 77.2500 192.9000 78.7500 ;
	    RECT 167.1000 77.1000 168.9000 77.2500 ;
	    RECT 191.1000 77.1000 192.9000 77.2500 ;
	    RECT 71.1000 72.7500 72.9000 72.9000 ;
	    RECT 80.7000 72.7500 82.5000 72.9000 ;
	    RECT 71.1000 71.2500 82.5000 72.7500 ;
	    RECT 71.1000 71.1000 72.9000 71.2500 ;
	    RECT 80.7000 71.1000 82.5000 71.2500 ;
	    RECT 95.1000 72.7500 96.9000 72.9000 ;
	    RECT 121.5000 72.7500 123.3000 72.9000 ;
	    RECT 95.1000 71.2500 123.3000 72.7500 ;
	    RECT 95.1000 71.1000 96.9000 71.2500 ;
	    RECT 121.5000 71.1000 123.3000 71.2500 ;
	    RECT 147.9000 72.7500 149.7000 72.9000 ;
	    RECT 155.1000 72.7500 156.9000 72.9000 ;
	    RECT 147.9000 71.2500 156.9000 72.7500 ;
	    RECT 147.9000 71.1000 149.7000 71.2500 ;
	    RECT 155.1000 71.1000 156.9000 71.2500 ;
	    RECT 140.7000 66.7500 142.5000 66.9000 ;
	    RECT 152.7000 66.7500 154.5000 66.9000 ;
	    RECT 162.3000 66.7500 164.1000 66.9000 ;
	    RECT 140.7000 65.2500 164.1000 66.7500 ;
	    RECT 140.7000 65.1000 142.5000 65.2500 ;
	    RECT 152.7000 65.1000 154.5000 65.2500 ;
	    RECT 162.3000 65.1000 164.1000 65.2500 ;
	    RECT 51.6000 60.6000 58.8000 62.4000 ;
	    RECT 126.3000 60.7500 128.1000 60.9000 ;
	    RECT 143.1000 60.7500 144.9000 60.9000 ;
	    RECT 126.3000 59.2500 144.9000 60.7500 ;
	    RECT 126.3000 59.1000 128.1000 59.2500 ;
	    RECT 143.1000 59.1000 144.9000 59.2500 ;
	    RECT 104.7000 54.7500 106.5000 54.9000 ;
	    RECT 109.5000 54.7500 111.3000 54.9000 ;
	    RECT 104.7000 53.2500 111.3000 54.7500 ;
	    RECT 104.7000 53.1000 106.5000 53.2500 ;
	    RECT 109.5000 53.1000 111.3000 53.2500 ;
	    RECT 150.3000 54.7500 152.1000 54.9000 ;
	    RECT 159.9000 54.7500 161.7000 54.9000 ;
	    RECT 150.3000 53.2500 161.7000 54.7500 ;
	    RECT 150.3000 53.1000 152.1000 53.2500 ;
	    RECT 159.9000 53.1000 161.7000 53.2500 ;
	    RECT 23.1000 48.7500 24.9000 48.9000 ;
	    RECT 32.7000 48.7500 34.5000 48.9000 ;
	    RECT 23.1000 47.2500 34.5000 48.7500 ;
	    RECT 23.1000 47.1000 24.9000 47.2500 ;
	    RECT 32.7000 47.1000 34.5000 47.2500 ;
	    RECT 39.9000 48.7500 41.7000 48.9000 ;
	    RECT 49.5000 48.7500 51.3000 48.9000 ;
	    RECT 39.9000 47.2500 51.3000 48.7500 ;
	    RECT 39.9000 47.1000 41.7000 47.2500 ;
	    RECT 49.5000 47.1000 51.3000 47.2500 ;
	    RECT 61.5000 48.7500 63.3000 48.9000 ;
	    RECT 71.1000 48.7500 72.9000 48.9000 ;
	    RECT 61.5000 47.2500 72.9000 48.7500 ;
	    RECT 61.5000 47.1000 63.3000 47.2500 ;
	    RECT 71.1000 47.1000 72.9000 47.2500 ;
	    RECT 75.9000 48.7500 77.7000 48.9000 ;
	    RECT 80.7000 48.7500 82.5000 48.9000 ;
	    RECT 85.5000 48.7500 87.3000 48.9000 ;
	    RECT 75.9000 47.2500 87.3000 48.7500 ;
	    RECT 75.9000 47.1000 77.7000 47.2500 ;
	    RECT 80.7000 47.1000 82.5000 47.2500 ;
	    RECT 85.5000 47.1000 87.3000 47.2500 ;
	    RECT 97.5000 48.7500 99.3000 48.9000 ;
	    RECT 102.3000 48.7500 104.1000 48.9000 ;
	    RECT 97.5000 47.2500 104.1000 48.7500 ;
	    RECT 97.5000 47.1000 99.3000 47.2500 ;
	    RECT 102.3000 47.1000 104.1000 47.2500 ;
	    RECT 109.5000 48.7500 111.3000 48.9000 ;
	    RECT 123.9000 48.7500 125.7000 48.9000 ;
	    RECT 147.9000 48.7500 149.7000 48.9000 ;
	    RECT 176.7000 48.7500 178.5000 48.9000 ;
	    RECT 109.5000 47.2500 178.5000 48.7500 ;
	    RECT 109.5000 47.1000 111.3000 47.2500 ;
	    RECT 123.9000 47.1000 125.7000 47.2500 ;
	    RECT 147.9000 47.1000 149.7000 47.2500 ;
	    RECT 176.7000 47.1000 178.5000 47.2500 ;
	    RECT 8.7000 44.1000 10.5000 45.9000 ;
	    RECT 171.9000 44.1000 173.7000 45.9000 ;
	    RECT 8.8500 42.7500 10.3500 44.1000 ;
	    RECT 25.5000 42.7500 27.3000 42.9000 ;
	    RECT 8.8500 41.2500 27.3000 42.7500 ;
	    RECT 25.5000 41.1000 27.3000 41.2500 ;
	    RECT 42.3000 42.7500 44.1000 42.9000 ;
	    RECT 78.3000 42.7500 80.1000 42.9000 ;
	    RECT 42.3000 41.2500 80.1000 42.7500 ;
	    RECT 42.3000 41.1000 44.1000 41.2500 ;
	    RECT 78.3000 41.1000 80.1000 41.2500 ;
	    RECT 92.7000 42.7500 94.5000 42.9000 ;
	    RECT 97.5000 42.7500 99.3000 42.9000 ;
	    RECT 92.7000 41.2500 99.3000 42.7500 ;
	    RECT 92.7000 41.1000 94.5000 41.2500 ;
	    RECT 97.5000 41.1000 99.3000 41.2500 ;
	    RECT 102.3000 42.7500 104.1000 42.9000 ;
	    RECT 111.9000 42.7500 113.7000 42.9000 ;
	    RECT 102.3000 41.2500 113.7000 42.7500 ;
	    RECT 102.3000 41.1000 104.1000 41.2500 ;
	    RECT 111.9000 41.1000 113.7000 41.2500 ;
	    RECT 119.1000 42.7500 120.9000 42.9000 ;
	    RECT 128.7000 42.7500 130.5000 42.9000 ;
	    RECT 119.1000 41.2500 130.5000 42.7500 ;
	    RECT 119.1000 41.1000 120.9000 41.2500 ;
	    RECT 128.7000 41.1000 130.5000 41.2500 ;
	    RECT 143.1000 42.7500 144.9000 42.9000 ;
	    RECT 150.3000 42.7500 152.1000 42.9000 ;
	    RECT 143.1000 41.2500 152.1000 42.7500 ;
	    RECT 172.0500 42.7500 173.5500 44.1000 ;
	    RECT 183.9000 42.7500 185.7000 42.9000 ;
	    RECT 172.0500 41.2500 185.7000 42.7500 ;
	    RECT 143.1000 41.1000 144.9000 41.2500 ;
	    RECT 150.3000 41.1000 152.1000 41.2500 ;
	    RECT 183.9000 41.1000 185.7000 41.2500 ;
	    RECT 75.9000 36.7500 77.7000 36.9000 ;
	    RECT 80.7000 36.7500 82.5000 36.9000 ;
	    RECT 75.9000 35.2500 82.5000 36.7500 ;
	    RECT 75.9000 35.1000 77.7000 35.2500 ;
	    RECT 80.7000 35.1000 82.5000 35.2500 ;
	    RECT 114.3000 36.7500 116.1000 36.9000 ;
	    RECT 126.3000 36.7500 128.1000 36.9000 ;
	    RECT 114.3000 35.2500 128.1000 36.7500 ;
	    RECT 114.3000 35.1000 116.1000 35.2500 ;
	    RECT 126.3000 35.1000 128.1000 35.2500 ;
	    RECT 157.5000 36.7500 159.3000 36.9000 ;
	    RECT 167.1000 36.7500 168.9000 36.9000 ;
	    RECT 157.5000 35.2500 168.9000 36.7500 ;
	    RECT 157.5000 35.1000 159.3000 35.2500 ;
	    RECT 167.1000 35.1000 168.9000 35.2500 ;
	    RECT 66.3000 30.7500 68.1000 30.9000 ;
	    RECT 71.1000 30.7500 72.9000 30.9000 ;
	    RECT 95.1000 30.7500 96.9000 30.9000 ;
	    RECT 66.3000 29.2500 96.9000 30.7500 ;
	    RECT 133.2000 30.6000 140.4000 32.4000 ;
	    RECT 181.5000 30.7500 183.3000 30.9000 ;
	    RECT 186.3000 30.7500 188.1000 30.9000 ;
	    RECT 66.3000 29.1000 68.1000 29.2500 ;
	    RECT 71.1000 29.1000 72.9000 29.2500 ;
	    RECT 95.1000 29.1000 96.9000 29.2500 ;
	    RECT 181.5000 29.2500 188.1000 30.7500 ;
	    RECT 181.5000 29.1000 183.3000 29.2500 ;
	    RECT 186.3000 29.1000 188.1000 29.2500 ;
	    RECT 3.9000 24.7500 5.7000 24.9000 ;
	    RECT 15.9000 24.7500 17.7000 24.9000 ;
	    RECT 3.9000 23.2500 17.7000 24.7500 ;
	    RECT 3.9000 23.1000 5.7000 23.2500 ;
	    RECT 15.9000 23.1000 17.7000 23.2500 ;
	    RECT 20.7000 24.7500 22.5000 24.9000 ;
	    RECT 25.5000 24.7500 27.3000 24.9000 ;
	    RECT 20.7000 23.2500 27.3000 24.7500 ;
	    RECT 20.7000 23.1000 22.5000 23.2500 ;
	    RECT 25.5000 23.1000 27.3000 23.2500 ;
	    RECT 32.7000 24.7500 34.5000 24.9000 ;
	    RECT 44.7000 24.7500 46.5000 24.9000 ;
	    RECT 32.7000 23.2500 46.5000 24.7500 ;
	    RECT 32.7000 23.1000 34.5000 23.2500 ;
	    RECT 44.7000 23.1000 46.5000 23.2500 ;
	    RECT 54.3000 24.7500 56.1000 24.9000 ;
	    RECT 78.3000 24.7500 80.1000 24.9000 ;
	    RECT 54.3000 23.2500 80.1000 24.7500 ;
	    RECT 54.3000 23.1000 56.1000 23.2500 ;
	    RECT 78.3000 23.1000 80.1000 23.2500 ;
	    RECT 140.7000 24.7500 142.5000 24.9000 ;
	    RECT 152.7000 24.7500 154.5000 24.9000 ;
	    RECT 159.9000 24.7500 161.7000 24.9000 ;
	    RECT 140.7000 23.2500 161.7000 24.7500 ;
	    RECT 140.7000 23.1000 142.5000 23.2500 ;
	    RECT 152.7000 23.1000 154.5000 23.2500 ;
	    RECT 159.9000 23.1000 161.7000 23.2500 ;
	    RECT 11.1000 18.7500 12.9000 18.9000 ;
	    RECT 15.9000 18.7500 17.7000 18.9000 ;
	    RECT 11.1000 17.2500 17.7000 18.7500 ;
	    RECT 11.1000 17.1000 12.9000 17.2500 ;
	    RECT 15.9000 17.1000 17.7000 17.2500 ;
	    RECT 20.7000 18.7500 22.5000 18.9000 ;
	    RECT 37.5000 18.7500 39.3000 18.9000 ;
	    RECT 56.7000 18.7500 58.5000 18.9000 ;
	    RECT 20.7000 17.2500 58.5000 18.7500 ;
	    RECT 20.7000 17.1000 22.5000 17.2500 ;
	    RECT 37.5000 17.1000 39.3000 17.2500 ;
	    RECT 56.7000 17.1000 58.5000 17.2500 ;
	    RECT 138.3000 18.7500 140.1000 18.9000 ;
	    RECT 143.1000 18.7500 144.9000 18.9000 ;
	    RECT 138.3000 17.2500 144.9000 18.7500 ;
	    RECT 138.3000 17.1000 140.1000 17.2500 ;
	    RECT 143.1000 17.1000 144.9000 17.2500 ;
	    RECT 147.9000 18.7500 149.7000 18.9000 ;
	    RECT 152.7000 18.7500 154.5000 18.9000 ;
	    RECT 147.9000 17.2500 154.5000 18.7500 ;
	    RECT 147.9000 17.1000 149.7000 17.2500 ;
	    RECT 152.7000 17.1000 154.5000 17.2500 ;
	    RECT 174.3000 12.7500 176.1000 12.9000 ;
	    RECT 179.1000 12.7500 180.9000 12.9000 ;
	    RECT 174.3000 11.2500 180.9000 12.7500 ;
	    RECT 174.3000 11.1000 176.1000 11.2500 ;
	    RECT 179.1000 11.1000 180.9000 11.2500 ;
	    RECT 51.6000 0.6000 58.8000 2.4000 ;
   END
END adder
