magic
tech scmos
timestamp 1590329367
<< metal1 >>
rect -2 97 26 103
rect 2 57 6 94
rect 10 60 14 94
rect 2 54 13 57
rect 18 54 22 94
rect 10 51 13 54
rect 10 47 16 51
rect 2 43 6 47
rect 2 39 6 40
rect 10 32 13 47
rect 19 43 22 54
rect 18 40 22 43
rect 18 33 22 37
rect 2 29 13 32
rect 2 6 6 29
rect 10 6 14 26
rect 18 6 22 30
rect -2 -3 26 3
<< labels >>
rlabel metal1 2 43 6 47 6 A
port 1 nsew default input
rlabel metal1 -2 -3 26 3 8 gnd
port 2 nsew ground bidirectional
rlabel metal1 18 33 22 37 6 Y
port 3 nsew default output
rlabel metal1 -2 97 26 103 6 vdd
port 4 nsew power bidirectional
<< properties >>
string LEFclass CORE
string LEFsite core
string LEFview TRUE
string FIXED_BBOX 0 0 24 100
string LEFsymmetry X Y
<< end >>
