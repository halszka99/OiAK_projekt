magic
tech scmos
timestamp 1590329367
<< metal1 >>
rect -2 97 58 103
rect 2 54 6 94
rect 10 54 14 94
rect 25 74 31 94
rect 18 53 22 57
rect 42 54 46 94
rect 2 49 6 50
rect 13 50 15 51
rect 13 47 22 50
rect 30 47 47 51
rect 50 50 54 94
rect 21 43 25 44
rect 50 43 54 47
rect 6 40 25 43
rect 6 33 7 37
rect 10 33 14 37
rect 29 36 33 41
rect 37 40 47 42
rect 37 38 54 40
rect 17 33 33 36
rect 2 6 6 26
rect 10 6 14 26
rect 22 23 26 33
rect 25 6 31 16
rect 42 6 46 26
rect 50 6 54 38
rect -2 -3 58 3
<< m2contact >>
rect 26 70 30 74
rect 2 50 6 54
rect 26 47 30 51
rect 2 40 6 44
rect 2 26 6 30
rect 26 16 30 20
<< metal2 >>
rect 2 44 6 50
rect 2 30 6 40
rect 26 51 30 70
rect 26 20 30 47
<< labels >>
rlabel metal1 50 43 54 47 6 Q
port 1 nsew default output
rlabel metal1 10 33 14 37 6 CLK
port 2 nsew default input
rlabel metal1 18 53 22 57 6 D
port 3 nsew default input
rlabel metal1 -2 -3 58 3 8 gnd
port 4 nsew ground bidirectional
rlabel metal1 -2 97 58 103 6 vdd
port 5 nsew power bidirectional
<< properties >>
string LEFclass CORE
string LEFsite core
string LEFview TRUE
string FIXED_BBOX 0 0 56 100
string LEFsymmetry X Y
<< end >>
