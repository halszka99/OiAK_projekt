magic
tech scmos
timestamp 1590329367
<< metal1 >>
rect -2 97 74 103
rect 2 54 6 94
rect 10 51 14 94
rect 18 54 22 94
rect 26 51 30 94
rect 34 54 38 94
rect 42 51 46 94
rect 50 54 54 94
rect 58 51 62 94
rect 66 54 70 94
rect 10 47 19 51
rect 26 47 37 51
rect 42 47 53 51
rect 58 50 70 51
rect 58 47 63 50
rect 15 40 19 47
rect 33 40 37 47
rect 49 40 53 47
rect 66 43 70 47
rect 2 33 6 37
rect 9 36 11 40
rect 15 36 28 40
rect 33 36 45 40
rect 49 36 62 40
rect 15 33 19 36
rect 33 33 37 36
rect 49 33 53 36
rect 66 33 70 40
rect 10 29 19 33
rect 26 29 37 33
rect 42 29 53 33
rect 58 29 70 33
rect 2 6 6 26
rect 10 6 14 29
rect 18 6 22 26
rect 26 6 30 29
rect 34 6 38 26
rect 42 6 46 29
rect 50 6 54 26
rect 58 6 62 29
rect 66 6 70 26
rect -2 -3 74 3
<< labels >>
rlabel metal1 2 33 6 37 6 A
port 1 nsew default input
rlabel metal1 -2 -3 74 3 8 gnd
port 2 nsew ground bidirectional
rlabel metal1 66 43 70 47 6 Y
port 3 nsew default output
rlabel metal1 -2 97 74 103 6 vdd
port 4 nsew power bidirectional
<< properties >>
string LEFclass CORE
string LEFsite core
string LEFview TRUE
string FIXED_BBOX 0 0 72 100
string LEFsymmetry X Y
<< end >>
