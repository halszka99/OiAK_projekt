magic
tech scmos
timestamp 1590329367
<< metal1 >>
rect -2 97 26 103
rect 2 54 6 94
rect 15 58 19 94
rect 10 54 19 58
rect 11 40 14 54
rect 18 50 22 51
rect 18 43 22 47
rect 10 33 14 37
rect 2 23 6 27
rect 2 19 6 20
rect 11 16 14 30
rect 2 6 6 16
rect 10 6 14 16
rect 18 6 22 16
rect -2 -3 26 3
<< labels >>
rlabel metal1 2 23 6 27 6 A
port 1 nsew default input
rlabel metal1 18 43 22 47 6 B
port 2 nsew default input
rlabel metal1 -2 -3 26 3 8 gnd
port 3 nsew ground bidirectional
rlabel metal1 10 33 14 37 6 Y
port 4 nsew default output
rlabel metal1 -2 97 26 103 6 vdd
port 5 nsew power bidirectional
<< properties >>
string LEFclass CORE
string LEFsite core
string LEFview TRUE
string FIXED_BBOX 0 0 24 100
string LEFsymmetry X Y
<< end >>
