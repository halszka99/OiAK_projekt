magic
tech scmos
timestamp 1590329367
<< metal1 >>
rect -2 97 34 103
rect 2 54 6 94
rect 15 57 19 94
rect 23 74 27 94
rect 22 63 26 67
rect 23 60 26 63
rect 15 54 20 57
rect 10 43 14 47
rect 10 39 14 40
rect 17 37 20 54
rect 26 53 30 57
rect 2 33 6 37
rect 9 31 10 36
rect 17 33 23 37
rect 26 33 30 37
rect 3 26 21 28
rect 26 26 29 30
rect 2 25 22 26
rect 2 6 6 25
rect 10 6 14 22
rect 18 6 22 25
rect 26 6 30 26
rect -2 -3 34 3
<< labels >>
rlabel metal1 2 33 6 37 6 A
port 1 nsew default input
rlabel metal1 10 43 14 47 6 B
port 2 nsew default input
rlabel metal1 26 53 30 57 6 C
port 3 nsew default input
rlabel metal1 -2 -3 34 3 8 gnd
port 4 nsew ground bidirectional
rlabel metal1 26 33 30 37 6 Y
port 5 nsew default output
rlabel metal1 -2 97 34 103 6 vdd
port 6 nsew power bidirectional
<< properties >>
string LEFclass CORE
string LEFsite core
string LEFview TRUE
string FIXED_BBOX 0 0 32 100
string LEFsymmetry X Y
<< end >>
