VERSION 5.3 ;
   NAMESCASESENSITIVE ON ;
   NOWIREEXTENSIONATPIN ON ;
   DIVIDERCHAR "/" ;
   BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO dot
   CLASS BLOCK ;
   FOREIGN dot ;
   ORIGIN 3.1500 -0.6000 ;
   SIZE 66.3000 BY 42.0000 ;
   PIN Gh
      PORT
         LAYER metal1 ;
	    RECT 42.6000 42.4500 43.8000 42.6000 ;
	    RECT 49.8000 42.4500 51.0000 42.6000 ;
	    RECT 42.6000 41.5500 51.0000 42.4500 ;
	    RECT 42.6000 41.4000 43.8000 41.5500 ;
	    RECT 49.8000 41.4000 51.0000 41.5500 ;
	    RECT 49.8000 23.4000 51.0000 24.6000 ;
         LAYER metal2 ;
	    RECT 42.6000 41.4000 43.8000 42.6000 ;
	    RECT 49.8000 41.4000 51.0000 42.6000 ;
	    RECT 42.7500 35.5500 43.6500 41.4000 ;
	    RECT 49.9500 24.6000 50.8500 41.4000 ;
	    RECT 49.8000 23.4000 51.0000 24.6000 ;
      END
   END Gh
   PIN Ph
      PORT
         LAYER metal1 ;
	    RECT 23.4000 20.4000 24.6000 21.6000 ;
	    RECT 23.4000 15.4500 24.6000 15.6000 ;
	    RECT 25.8000 15.4500 27.0000 15.6000 ;
	    RECT 23.4000 14.5500 27.0000 15.4500 ;
	    RECT 23.4000 14.4000 24.6000 14.5500 ;
	    RECT 25.8000 14.4000 27.0000 14.5500 ;
         LAYER metal2 ;
	    RECT 16.3500 24.6000 17.2500 36.4500 ;
	    RECT 16.2000 23.4000 17.4000 24.6000 ;
	    RECT 23.4000 23.4000 24.6000 24.6000 ;
	    RECT 23.5500 21.6000 24.4500 23.4000 ;
	    RECT 23.4000 20.4000 24.6000 21.6000 ;
	    RECT 23.5500 15.6000 24.4500 20.4000 ;
	    RECT 23.4000 14.4000 24.6000 15.6000 ;
         LAYER metal3 ;
	    RECT 15.9000 24.7500 17.7000 24.9000 ;
	    RECT 23.1000 24.7500 24.9000 24.9000 ;
	    RECT 15.9000 23.2500 24.9000 24.7500 ;
	    RECT 15.9000 23.1000 17.7000 23.2500 ;
	    RECT 23.1000 23.1000 24.9000 23.2500 ;
      END
   END Ph
   PIN Gl
      PORT
         LAYER metal1 ;
	    RECT 30.6000 20.4000 31.8000 21.6000 ;
         LAYER metal2 ;
	    RECT 30.7500 21.6000 31.6500 36.4500 ;
	    RECT 30.6000 20.4000 31.8000 21.6000 ;
      END
   END Gl
   PIN Pl
      PORT
         LAYER metal1 ;
	    RECT 21.0000 17.4000 22.2000 18.6000 ;
         LAYER metal2 ;
	    RECT 21.0000 17.4000 22.2000 18.6000 ;
	    RECT 21.1500 12.6000 22.0500 17.4000 ;
	    RECT 21.0000 11.4000 22.2000 12.6000 ;
         LAYER metal3 ;
	    RECT -3.1500 12.7500 -1.6500 18.7500 ;
	    RECT 20.7000 12.7500 22.5000 12.9000 ;
	    RECT -3.1500 11.2500 22.5000 12.7500 ;
	    RECT 20.7000 11.1000 22.5000 11.2500 ;
      END
   END Pl
   PIN Ghl
      PORT
         LAYER metal1 ;
	    RECT 57.0000 20.4000 58.2000 21.6000 ;
         LAYER metal2 ;
	    RECT 57.0000 20.4000 58.2000 21.6000 ;
	    RECT 57.1500 18.6000 58.0500 20.4000 ;
	    RECT 57.0000 17.4000 58.2000 18.6000 ;
         LAYER metal3 ;
	    RECT 56.7000 18.7500 58.5000 18.9000 ;
	    RECT 61.6500 18.7500 63.1500 24.7500 ;
	    RECT 56.7000 17.2500 63.1500 18.7500 ;
	    RECT 56.7000 17.1000 58.5000 17.2500 ;
      END
   END Ghl
   PIN Phl
      PORT
         LAYER metal1 ;
	    RECT 1.8000 20.4000 3.0000 21.6000 ;
         LAYER metal2 ;
	    RECT 1.8000 29.4000 3.0000 30.6000 ;
	    RECT 1.9500 21.6000 2.8500 29.4000 ;
	    RECT 1.8000 20.4000 3.0000 21.6000 ;
         LAYER metal3 ;
	    RECT 1.5000 30.7500 3.3000 30.9000 ;
	    RECT -3.1500 29.2500 3.3000 30.7500 ;
	    RECT -3.1500 23.2500 -1.6500 29.2500 ;
	    RECT 1.5000 29.1000 3.3000 29.2500 ;
      END
   END Phl
   OBS
         LAYER metal1 ;
	    RECT 0.6000 30.6000 59.4000 32.4000 ;
	    RECT 1.8000 22.5000 3.0000 29.7000 ;
	    RECT 4.2000 23.7000 5.4000 29.7000 ;
	    RECT 6.6000 22.8000 7.8000 29.7000 ;
	    RECT 17.1000 25.2000 18.3000 29.7000 ;
	    RECT 4.5000 21.9000 7.8000 22.8000 ;
	    RECT 16.2000 23.7000 18.3000 25.2000 ;
	    RECT 19.5000 24.0000 20.7000 29.7000 ;
	    RECT 23.4000 23.7000 24.6000 29.7000 ;
	    RECT 26.7000 24.6000 27.9000 29.7000 ;
	    RECT 26.7000 23.7000 29.4000 24.6000 ;
	    RECT 30.6000 23.7000 31.8000 29.7000 ;
	    RECT 33.9000 24.6000 35.1000 29.7000 ;
	    RECT 33.9000 23.7000 36.6000 24.6000 ;
	    RECT 37.8000 23.7000 39.0000 29.7000 ;
	    RECT 1.8000 18.6000 3.0000 19.5000 ;
	    RECT 1.8000 15.3000 2.7000 18.6000 ;
	    RECT 4.5000 17.4000 5.4000 21.9000 ;
	    RECT 6.6000 19.5000 7.8000 19.8000 ;
	    RECT 16.2000 19.5000 17.1000 23.7000 ;
	    RECT 23.4000 23.4000 24.3000 23.7000 ;
	    RECT 21.6000 22.8000 24.3000 23.4000 ;
	    RECT 18.0000 22.5000 24.3000 22.8000 ;
	    RECT 18.0000 21.9000 22.5000 22.5000 ;
	    RECT 18.0000 21.6000 19.2000 21.9000 ;
	    RECT 6.6000 18.4500 7.8000 18.6000 ;
	    RECT 16.2000 18.4500 17.4000 18.6000 ;
	    RECT 6.6000 17.5500 17.4000 18.4500 ;
	    RECT 6.6000 17.4000 7.8000 17.5500 ;
	    RECT 16.2000 17.4000 17.4000 17.5500 ;
	    RECT 3.6000 16.2000 5.4000 17.4000 ;
	    RECT 18.3000 16.5000 19.2000 21.6000 ;
	    RECT 20.4000 20.7000 21.6000 21.0000 ;
	    RECT 20.4000 19.8000 21.9000 20.7000 ;
	    RECT 21.0000 19.5000 21.9000 19.8000 ;
	    RECT 28.2000 19.5000 29.4000 23.7000 ;
	    RECT 30.6000 22.5000 31.8000 22.8000 ;
	    RECT 35.4000 19.5000 36.6000 23.7000 ;
	    RECT 37.8000 22.5000 39.0000 22.8000 ;
	    RECT 47.4000 22.5000 48.6000 29.7000 ;
	    RECT 49.8000 26.7000 51.0000 29.7000 ;
	    RECT 49.8000 25.5000 51.0000 25.8000 ;
	    RECT 52.2000 22.8000 53.4000 29.7000 ;
	    RECT 54.6000 23.7000 55.8000 29.7000 ;
	    RECT 52.2000 21.9000 55.5000 22.8000 ;
	    RECT 57.0000 22.5000 58.2000 29.7000 ;
	    RECT 37.8000 21.4500 39.0000 21.6000 ;
	    RECT 47.4000 21.4500 48.6000 21.6000 ;
	    RECT 37.8000 20.5500 48.6000 21.4500 ;
	    RECT 37.8000 20.4000 39.0000 20.5500 ;
	    RECT 47.4000 20.4000 48.6000 20.5500 ;
	    RECT 52.2000 19.5000 53.4000 19.8000 ;
	    RECT 23.4000 19.2000 24.6000 19.5000 ;
	    RECT 28.2000 18.4500 29.4000 18.6000 ;
	    RECT 35.4000 18.4500 36.6000 18.6000 ;
	    RECT 45.0000 18.4500 46.2000 18.6000 ;
	    RECT 28.2000 17.5500 34.0500 18.4500 ;
	    RECT 28.2000 17.4000 29.4000 17.5500 ;
	    RECT 4.5000 15.3000 5.4000 16.2000 ;
	    RECT 16.2000 15.3000 17.1000 16.5000 ;
	    RECT 18.3000 15.6000 21.9000 16.5000 ;
	    RECT 1.8000 3.3000 3.0000 15.3000 ;
	    RECT 4.5000 14.4000 7.8000 15.3000 ;
	    RECT 4.2000 3.3000 5.4000 13.5000 ;
	    RECT 6.6000 3.3000 7.8000 14.4000 ;
	    RECT 16.2000 3.3000 17.4000 15.3000 ;
	    RECT 18.6000 3.3000 19.8000 14.7000 ;
	    RECT 21.0000 9.3000 21.9000 15.6000 ;
	    RECT 25.8000 13.2000 27.0000 13.5000 ;
	    RECT 21.0000 3.3000 22.2000 9.3000 ;
	    RECT 23.4000 3.3000 24.6000 9.3000 ;
	    RECT 25.8000 3.3000 27.0000 9.3000 ;
	    RECT 28.2000 3.3000 29.4000 16.5000 ;
	    RECT 33.1500 15.6000 34.0500 17.5500 ;
	    RECT 35.4000 17.5500 46.2000 18.4500 ;
	    RECT 35.4000 17.4000 36.6000 17.5500 ;
	    RECT 45.0000 17.4000 46.2000 17.5500 ;
	    RECT 33.0000 14.4000 34.2000 15.6000 ;
	    RECT 33.0000 13.2000 34.2000 13.5000 ;
	    RECT 30.6000 3.3000 31.8000 9.3000 ;
	    RECT 33.0000 3.3000 34.2000 9.3000 ;
	    RECT 35.4000 3.3000 36.6000 16.5000 ;
	    RECT 37.8000 3.3000 39.0000 9.3000 ;
	    RECT 47.4000 3.3000 48.6000 19.5000 ;
	    RECT 52.2000 17.4000 53.4000 18.6000 ;
	    RECT 54.6000 17.4000 55.5000 21.9000 ;
	    RECT 57.0000 18.6000 58.2000 19.5000 ;
	    RECT 54.6000 16.2000 56.4000 17.4000 ;
	    RECT 54.6000 15.3000 55.5000 16.2000 ;
	    RECT 57.3000 15.3000 58.2000 18.6000 ;
	    RECT 52.2000 14.4000 55.5000 15.3000 ;
	    RECT 49.8000 3.3000 51.0000 9.3000 ;
	    RECT 52.2000 3.3000 53.4000 14.4000 ;
	    RECT 54.6000 3.3000 55.8000 13.5000 ;
	    RECT 57.0000 3.3000 58.2000 15.3000 ;
	    RECT 0.6000 0.6000 59.4000 2.4000 ;
         LAYER metal2 ;
	    RECT 39.6000 30.6000 46.8000 32.4000 ;
	    RECT 45.0000 17.4000 46.2000 18.6000 ;
	    RECT 52.2000 17.4000 53.4000 18.6000 ;
	    RECT 8.4000 0.6000 15.6000 2.4000 ;
         LAYER metal3 ;
	    RECT 39.6000 30.6000 46.8000 32.4000 ;
	    RECT 44.7000 18.7500 46.5000 18.9000 ;
	    RECT 51.9000 18.7500 53.7000 18.9000 ;
	    RECT 44.7000 17.2500 53.7000 18.7500 ;
	    RECT 44.7000 17.1000 46.5000 17.2500 ;
	    RECT 51.9000 17.1000 53.7000 17.2500 ;
	    RECT 8.4000 0.6000 15.6000 2.4000 ;
   END
END dot
