magic
tech scmos
timestamp 1590329367
<< metal1 >>
rect -2 97 66 103
rect 2 64 6 94
rect 10 64 14 94
rect 18 91 38 94
rect 18 64 22 91
rect 26 64 30 88
rect 34 65 38 91
rect 43 91 61 94
rect 43 90 46 91
rect 3 61 6 64
rect 18 61 21 64
rect 3 58 21 61
rect 27 62 30 64
rect 42 62 46 90
rect 58 90 61 91
rect 27 60 46 62
rect 50 60 54 88
rect 58 60 62 90
rect 27 59 45 60
rect 37 53 47 56
rect 50 53 54 57
rect 26 43 30 47
rect 33 43 34 47
rect 18 33 22 37
rect 25 33 26 37
rect 10 23 14 27
rect 17 23 19 27
rect 37 20 40 53
rect 20 17 40 20
rect 20 16 23 17
rect 10 6 14 16
rect 18 13 23 16
rect 34 16 40 17
rect 18 6 22 13
rect 26 6 30 14
rect 34 6 38 16
rect -2 -3 66 3
<< labels >>
rlabel metal1 10 23 14 27 6 A
port 1 nsew default input
rlabel metal1 18 33 22 37 6 B
port 2 nsew default input
rlabel metal1 26 43 30 47 6 C
port 3 nsew default input
rlabel metal1 -2 -3 66 3 8 gnd
port 4 nsew ground bidirectional
rlabel metal1 50 53 54 57 6 Y
port 5 nsew default output
rlabel metal1 -2 97 66 103 6 vdd
port 6 nsew power bidirectional
<< properties >>
string LEFclass CORE
string LEFsite core
string LEFview TRUE
string FIXED_BBOX 0 0 64 100
string LEFsymmetry X Y
<< end >>
