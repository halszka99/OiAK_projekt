magic
tech scmos
timestamp 1590329367
<< metal1 >>
rect -2 97 34 103
rect 2 74 6 94
rect 10 74 14 94
rect 18 74 22 94
rect 26 74 30 94
rect 11 71 14 74
rect 11 68 23 71
rect 27 70 30 74
rect 10 53 14 57
rect 13 49 17 50
rect 2 40 6 41
rect 2 33 6 37
rect 20 33 23 68
rect 26 63 30 67
rect 9 30 24 33
rect 9 29 12 30
rect 20 29 24 30
rect 3 26 12 29
rect 2 6 6 26
rect 15 6 19 26
rect 27 19 30 60
rect 23 16 30 19
rect 23 6 27 16
rect -2 -3 34 3
<< labels >>
rlabel metal1 2 33 6 37 6 A
port 1 nsew default input
rlabel metal1 10 53 14 57 6 B
port 2 nsew default input
rlabel metal1 -2 -3 34 3 8 gnd
port 3 nsew ground bidirectional
rlabel metal1 26 63 30 67 6 Y
port 4 nsew default output
rlabel metal1 -2 97 34 103 6 vdd
port 5 nsew power bidirectional
<< properties >>
string LEFclass CORE
string LEFsite core
string LEFview TRUE
string FIXED_BBOX 0 0 32 100
string LEFsymmetry X Y
<< end >>
