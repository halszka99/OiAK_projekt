magic
tech scmos
timestamp 1590329367
<< metal1 >>
rect -2 97 34 103
rect 2 74 6 94
rect 10 74 14 94
rect 11 53 14 74
rect 18 56 22 94
rect 26 54 30 94
rect 11 50 23 53
rect 27 50 30 54
rect 10 43 14 47
rect 2 40 6 41
rect 11 39 14 40
rect 2 33 6 37
rect 11 36 16 39
rect 12 35 16 36
rect 20 33 23 50
rect 26 43 30 47
rect 20 32 24 33
rect 9 30 24 32
rect 3 29 24 30
rect 3 27 12 29
rect 3 26 6 27
rect 27 26 30 40
rect 2 6 6 26
rect 15 6 19 25
rect 23 21 30 26
rect 23 6 27 21
rect -2 -3 34 3
<< labels >>
rlabel metal1 2 33 6 37 6 A
port 1 nsew default input
rlabel metal1 10 43 14 47 6 B
port 2 nsew default input
rlabel metal1 -2 -3 34 3 8 gnd
port 3 nsew ground bidirectional
rlabel metal1 26 43 30 47 6 Y
port 4 nsew default output
rlabel metal1 -2 97 34 103 6 vdd
port 5 nsew power bidirectional
<< properties >>
string LEFclass CORE
string LEFsite core
string LEFview TRUE
string FIXED_BBOX 0 0 32 100
string LEFsymmetry X Y
<< end >>
