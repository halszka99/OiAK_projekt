magic
tech scmos
timestamp 1590329367
<< metal1 >>
rect -2 97 58 103
rect 2 54 6 94
rect 10 54 14 94
rect 18 91 38 94
rect 18 54 22 91
rect 26 54 30 88
rect 34 58 38 91
rect 42 61 46 94
rect 50 58 54 94
rect 34 54 54 58
rect 2 50 6 51
rect 2 43 6 47
rect 10 45 13 54
rect 26 50 29 54
rect 10 41 14 45
rect 26 43 30 47
rect 2 33 5 40
rect 2 29 7 33
rect 10 26 13 41
rect 26 26 29 40
rect 45 33 47 37
rect 50 33 54 37
rect 34 26 54 29
rect 2 6 6 26
rect 10 6 14 26
rect 18 9 22 26
rect 26 12 30 26
rect 34 9 38 26
rect 51 23 54 26
rect 18 6 38 9
rect 42 6 46 23
rect 50 6 54 23
rect -2 -3 58 3
<< labels >>
rlabel metal1 50 33 54 37 6 A
port 1 nsew default input
rlabel metal1 2 43 6 47 6 EN
port 2 nsew default input
rlabel metal1 -2 -3 58 3 8 gnd
port 3 nsew ground bidirectional
rlabel metal1 26 43 30 47 6 Y
port 4 nsew default output
rlabel metal1 -2 97 58 103 6 vdd
port 5 nsew power bidirectional
<< properties >>
string LEFclass CORE
string LEFsite core
string LEFview TRUE
string FIXED_BBOX 0 0 56 100
string LEFsymmetry X Y
<< end >>
